********************************************
* Ansys RedHawk-SC Chip Power Model [ Ver 2.00 ]
* Generated at Mar 09 03:28:04 2024
* Version: 2021 R1.RD  RHEL6 (Sep 29 00:01:22 2020)
* Run directory:  /fs/mm_imp46/user/kuma/03_240203_wDFT_for_STAPI/flat2020R32_CLK2/gp/asim_power_scratch.gv_rmv.4803 
* CPM Options:  
* perform powermodel -nx 3 -ny 4 -no_afs -noglobal_gnd -pincurrent -emi -plocnames 
* Copyright (c) 2002-2020 ANSYS, Inc.
* Presimulation time  0.000000ps
********************************************


* Partitioning of flip chip bump pad area - Die Top View
* ------------------------------------
* | (0 Ny) | (1 Ny) | .... | (Nx Ny) |
* ------------------------------------
* | (0 ..) | (1 ..) | .... | (Nx ..) |
* ------------------------------------
* | (0  1) | (1  1) | .... | (Nx  1) |
* ------------------------------------
* | (0  0) | (1  0) | .... | (Nx  0) |
* ------------------------------------
* Begin Chip Package Protocol --->
 * generated by asim_power_model 

.subckt adsPowerModel_cpu
+ PAR_0_0_VDD075CPU PAR_1_0_VSS PAR_1_0_VDD075CPU PAR_2_0_VSS PAR_2_0_VDD075CPU 
+ PAR_0_1_VSS PAR_0_1_VDD075CPU PAR_1_1_VSS PAR_1_1_VDD075CPU PAR_2_1_VSS 
+ PAR_2_1_VDD075CPU PAR_0_2_VSS PAR_0_2_VDD075CPU PAR_1_2_VSS PAR_1_2_VDD075CPU 
+ PAR_2_2_VSS PAR_2_2_VDD075CPU PAR_0_3_VSS PAR_0_3_VDD075CPU PAR_1_3_VSS 
+ PAR_1_3_VDD075CPU PAR_0_0_VSS 

* No connection to global ground (Spice node 0) *
C0_1 PAR_0_0_VDD075CPU PAR_0_0_VSS 4.96053796593e-10
R_1_1 PAR_0_0_VDD075CPU n23 0.00130390726399
C_1_1 n23 PAR_0_0_VSS 1.35730155806e-08
R_2_1 PAR_0_0_VDD075CPU n24 0.00291206667173
C_2_1 n24 PAR_0_0_VSS 1.7469973393e-08
R_3_1 PAR_0_0_VDD075CPU n25 0.00195919055181
C_3_1 n25 PAR_0_0_VSS 4.97689573803e-08
R_4_1 PAR_0_0_VDD075CPU n26 0.633217809169
R_7_1 PAR_0_0_VDD075CPU n26 1688000
C_4_1 n26 PAR_0_0_VSS 3.81303525783e-10
R_5_1 PAR_0_0_VDD075CPU n27 2.78389763143
R_8_1 PAR_0_0_VDD075CPU n27 1778000
C_5_1 n27 PAR_0_0_VSS 3.61271928927e-10
R_6_1 PAR_0_0_VDD075CPU n28 27.4575065597
R_9_1 PAR_0_0_VDD075CPU n28 1889000
C_6_1 n28 PAR_0_0_VSS 1.99930614495e-10
G0_2 PAR_1_0_VSS PAR_0_0_VDD075CPU PAR_1_0_VSS PAR_0_0_VDD075CPU -2.15929114107
C0_2 PAR_1_0_VSS PAR_0_0_VDD075CPU 1.94819817883e-10
R_1_2 PAR_1_0_VSS n29 0.0389713812778
C_1_2 n29 PAR_0_0_VDD075CPU 4.98634888543e-10
R_2_2 PAR_1_0_VSS n30 0.113441747708
C_2_2 n30 PAR_0_0_VDD075CPU 5.66389527938e-10
R_3_2 PAR_1_0_VSS n31 0.0605333208254
C_3_2 n31 PAR_0_0_VDD075CPU 1.93856886381e-09
L_4_2 PAR_1_0_VSS n32 8.4222007075e-11
R_4_2 n32 PAR_0_0_VDD075CPU 0.478956075551
L_5_2 PAR_1_0_VSS n33 2.95490403732e-08
R_5_2 n33 PAR_0_0_VDD075CPU 16.0529286525
L_6_2 PAR_1_0_VSS n34 1.37130276903e-06
R_6_2 n34 PAR_0_0_VDD075CPU 109.612064237
R0_3 PAR_1_0_VSS PAR_0_0_VSS 0.00309801277074
R_1_3 PAR_1_0_VSS n35 0.0835978956757
C_1_3 n35 PAR_0_0_VSS 7.60618894085e-10
L_2_3 PAR_1_0_VSS n36 2.81472675652e-12
R_2_3 n36 PAR_0_0_VSS 0.0300270026145
R_3_3 PAR_1_0_VSS n37 0.0515873344
C_3_3 n37 PAR_0_0_VSS 3.38326535732e-09
L_4_3 PAR_1_0_VSS n38 1.0571862507e-10
R_4_3 n38 PAR_0_0_VSS 0.177479318888
L_5_3 PAR_1_0_VSS n39 1.06445740411e-09
R_5_3 n39 PAR_0_0_VSS 0.785745988494
R_6_3 PAR_1_0_VSS n40 6.67349628053
R_10_3 PAR_1_0_VSS n40 1666000
C_6_3 n40 PAR_0_0_VSS 1.5635426314e-09
R0_4 PAR_1_0_VDD075CPU PAR_0_0_VDD075CPU 0.00377083931658
C0_4 PAR_1_0_VDD075CPU PAR_0_0_VDD075CPU 5.61118462081e-11
L_1_4 PAR_1_0_VDD075CPU n41 4.26843747744e-13
R_1_4 n41 PAR_0_0_VDD075CPU 0.0252221904093
L_2_4 PAR_1_0_VDD075CPU n42 2.65877016186e-12
R_2_4 n42 PAR_0_0_VDD075CPU 0.0560136144529
L_3_4 PAR_1_0_VDD075CPU n43 3.41584319156e-12
R_3_4 n43 PAR_0_0_VDD075CPU 0.0327150507036
L_4_4 PAR_1_0_VDD075CPU n44 1.47072187487e-08
R_4_4 n44 PAR_0_0_VDD075CPU 32.0877397253
L_5_4 PAR_1_0_VDD075CPU n45 4.75696015681e-07
R_5_4 n45 PAR_0_0_VDD075CPU 237.974646806
L_6_4 PAR_1_0_VDD075CPU n46 5.57305619362e-05
R_6_4 n46 PAR_0_0_VDD075CPU 1702.44427048
G0_5 PAR_1_0_VDD075CPU PAR_1_0_VSS PAR_1_0_VDD075CPU PAR_1_0_VSS -0.0434495291161
C0_5 PAR_1_0_VDD075CPU PAR_1_0_VSS 1.29582666091e-09
R_1_5 PAR_1_0_VDD075CPU n47 0.0018914432404
C_1_5 n47 PAR_1_0_VSS 8.39525864326e-09
R_2_5 PAR_1_0_VDD075CPU n48 0.0033536931412
C_2_5 n48 PAR_1_0_VSS 1.57129373792e-08
R_3_5 PAR_1_0_VDD075CPU n49 0.00278965637502
C_3_5 n49 PAR_1_0_VSS 3.52231196821e-08
R_4_5 PAR_1_0_VDD075CPU n50 0.861196377161
C_4_5 n50 PAR_1_0_VSS 3.00337790385e-10
L_5_5 PAR_1_0_VDD075CPU n51 9.5734735734e-08
R_5_5 n51 PAR_1_0_VSS 23.0152078506
G0_6 PAR_1_0_VDD075CPU PAR_0_0_VSS PAR_1_0_VDD075CPU PAR_0_0_VSS -1.47959001681
C0_6 PAR_1_0_VDD075CPU PAR_0_0_VSS 3.02667489955e-10
R_1_6 PAR_1_0_VDD075CPU n52 0.00813901461702
C_1_6 n52 PAR_0_0_VSS 1.83031345522e-09
R_2_6 PAR_1_0_VDD075CPU n53 0.0449752661448
C_2_6 n53 PAR_0_0_VSS 1.1239568466e-09
R_3_6 PAR_1_0_VDD075CPU n54 0.0251607304292
C_3_6 n54 PAR_0_0_VSS 4.14725095142e-09
L_4_6 PAR_1_0_VDD075CPU n55 1.27315119803e-10
R_4_6 n55 PAR_0_0_VSS 0.675862899057
R_5_6 PAR_1_0_VDD075CPU n56 5.0120045578
C_5_6 n56 PAR_0_0_VSS 1.92083288234e-10
R_6_6 PAR_1_0_VDD075CPU n57 50.0826129531
C_6_6 n57 PAR_0_0_VSS 1.51481424901e-10
G0_7 PAR_2_0_VSS PAR_0_0_VDD075CPU PAR_2_0_VSS PAR_0_0_VDD075CPU -0.185935281097
C0_7 PAR_2_0_VSS PAR_0_0_VDD075CPU 2.44877549462e-10
R_1_7 PAR_2_0_VSS n58 2.4279039782
C_1_7 n58 PAR_0_0_VDD075CPU 4.47958871846e-11
R_2_7 PAR_2_0_VSS n59 3.3692378002
C_2_7 n59 PAR_0_0_VDD075CPU 1.81515720959e-10
L_3_7 PAR_2_0_VSS n60 8.25652814532e-09
R_3_7 n60 PAR_0_0_VDD075CPU 6.90008281729
L_4_7 PAR_2_0_VSS n61 9.37379545623e-08
R_4_7 n61 PAR_0_0_VDD075CPU 31.6024786943
L_5_7 PAR_2_0_VSS n62 1.41130382949e-06
R_5_7 n62 PAR_0_0_VDD075CPU 106.764613976
R0_8 PAR_2_0_VSS PAR_1_0_VSS 0.00378223518045
C0_8 PAR_2_0_VSS PAR_1_0_VSS 2.38856388885e-11
L_1_8 PAR_2_0_VSS n63 1.1094401385e-12
R_1_8 n63 PAR_1_0_VSS 0.0338691895787
L_2_8 PAR_2_0_VSS n64 3.02850676813e-12
R_2_8 n64 PAR_1_0_VSS 0.0321248424894
L_3_8 PAR_2_0_VSS n65 3.01138234038e-11
R_3_8 n65 PAR_1_0_VSS 0.131398832235
L_4_8 PAR_2_0_VSS n66 1.52198370337e-10
R_4_8 n66 PAR_1_0_VSS 0.18364947494
L_5_8 PAR_2_0_VSS n67 5.95458476255e-10
R_5_8 n67 PAR_1_0_VSS 0.354896418248
L_6_8 PAR_2_0_VSS n68 4.84390447541e-08
R_6_8 n68 PAR_1_0_VSS 4.60098372097
G0_9 PAR_2_0_VSS PAR_1_0_VDD075CPU PAR_2_0_VSS PAR_1_0_VDD075CPU -0.0951128229023
C0_9 PAR_2_0_VSS PAR_1_0_VDD075CPU 3.43912783647e-10
R_1_9 PAR_2_0_VSS n69 0.0214355261252
C_1_9 n69 PAR_1_0_VDD075CPU 1.49420098657e-09
R_2_9 PAR_2_0_VSS n70 0.0189676958283
C_2_9 n70 PAR_1_0_VDD075CPU 4.98514114182e-09
R_3_9 PAR_2_0_VSS n71 0.54419020717
C_3_9 n71 PAR_1_0_VDD075CPU 3.49131326205e-10
R_4_9 PAR_2_0_VSS n72 5.4589968732
C_4_9 n72 PAR_1_0_VDD075CPU 1.43985609705e-10
L_5_9 PAR_2_0_VSS n73 2.83059560199e-08
R_5_9 n73 PAR_1_0_VDD075CPU 10.513829186
R0_10 PAR_2_0_VSS PAR_0_0_VSS 2.88907907536
C0_10 PAR_2_0_VSS PAR_0_0_VSS 3.4542850749e-10
R_1_10 PAR_2_0_VSS n74 0.0220261664233
C_1_10 n74 PAR_0_0_VSS 8.63693503137e-10
R_2_10 PAR_2_0_VSS n75 0.154380184888
C_2_10 n75 PAR_0_0_VSS 4.26521150654e-10
R_3_10 PAR_2_0_VSS n76 0.172721248161
C_3_10 n76 PAR_0_0_VSS 1.28015683566e-09
R_4_10 PAR_2_0_VSS n77 0.0756764989001
C_4_10 n77 PAR_0_0_VSS 1.38003944812e-08
R_5_10 PAR_2_0_VSS n78 3.51348225761
C_5_10 n78 PAR_0_0_VSS 1.61323779104e-09
R_6_10 PAR_2_0_VSS n79 15.3306272776
C_6_10 n79 PAR_0_0_VSS 1.16723693388e-09
G0_11 PAR_2_0_VDD075CPU PAR_0_0_VDD075CPU PAR_2_0_VDD075CPU PAR_0_0_VDD075CPU -3.3666808249
C0_11 PAR_2_0_VDD075CPU PAR_0_0_VDD075CPU 1.49377590254e-10
R_1_11 PAR_2_0_VDD075CPU n80 0.554618150185
C_1_11 n80 PAR_0_0_VDD075CPU 4.5454773727e-11
L_2_11 PAR_2_0_VDD075CPU n81 4.50966142918e-11
R_2_11 n81 PAR_0_0_VDD075CPU 0.386595987771
R_3_11 PAR_2_0_VDD075CPU n82 0.734361339351
C_3_11 n82 PAR_0_0_VDD075CPU 3.56334794541e-10
L_4_11 PAR_2_0_VDD075CPU n83 9.03326326799e-10
R_4_11 n83 PAR_0_0_VDD075CPU 1.48055551025
R_5_11 PAR_2_0_VDD075CPU n84 4.95267618988
C_5_11 n84 PAR_0_0_VDD075CPU 6.56537002671e-10
L_6_11 PAR_2_0_VDD075CPU n85 8.19481919469e-08
R_6_11 n85 PAR_0_0_VDD075CPU 9.37601455519
G0_12 PAR_2_0_VDD075CPU PAR_1_0_VSS PAR_2_0_VDD075CPU PAR_1_0_VSS -0.626576726205
C0_12 PAR_2_0_VDD075CPU PAR_1_0_VSS 2.15126202549e-10
R_1_12 PAR_2_0_VDD075CPU n86 0.0449776646703
C_1_12 n86 PAR_1_0_VSS 4.71292952326e-10
R_2_12 PAR_2_0_VDD075CPU n87 0.0772166056442
C_2_12 n87 PAR_1_0_VSS 8.3682610166e-10
R_3_12 PAR_2_0_VDD075CPU n88 0.0542586183205
C_3_12 n88 PAR_1_0_VSS 2.08825392076e-09
L_4_12 PAR_2_0_VDD075CPU n89 4.03441249436e-10
R_4_12 n89 PAR_1_0_VSS 1.79855776959
L_5_12 PAR_2_0_VDD075CPU n90 3.21541407332e-08
R_5_12 n90 PAR_1_0_VSS 16.5055081628
L_6_12 PAR_2_0_VDD075CPU n91 1.37166163524e-06
R_6_12 n91 PAR_1_0_VSS 100.101623675
R0_13 PAR_2_0_VDD075CPU PAR_1_0_VDD075CPU 0.00375329317061
C0_13 PAR_2_0_VDD075CPU PAR_1_0_VDD075CPU 9.8193442637e-11
L_1_13 PAR_2_0_VDD075CPU n92 4.29167646748e-13
R_1_13 n92 PAR_1_0_VDD075CPU 0.0255217251869
L_2_13 PAR_2_0_VDD075CPU n93 2.54934331426e-12
R_2_13 n93 PAR_1_0_VDD075CPU 0.0505700496785
L_3_13 PAR_2_0_VDD075CPU n94 3.14136871479e-12
R_3_13 n94 PAR_1_0_VDD075CPU 0.0300384855622
L_4_13 PAR_2_0_VDD075CPU n95 7.4856998746e-09
R_4_13 n95 PAR_1_0_VDD075CPU 19.3058127814
L_5_13 PAR_2_0_VDD075CPU n96 1.45443642166e-07
R_5_13 n96 PAR_1_0_VDD075CPU 117.545691233
L_6_13 PAR_2_0_VDD075CPU n97 8.9546762945e-06
R_6_13 n97 PAR_1_0_VDD075CPU 800.701150717
G0_14 PAR_2_0_VDD075CPU PAR_2_0_VSS PAR_2_0_VDD075CPU PAR_2_0_VSS -0.057711649137
C0_14 PAR_2_0_VDD075CPU PAR_2_0_VSS 7.16883385448e-10
R_1_14 PAR_2_0_VDD075CPU n98 0.000956851202835
C_1_14 n98 PAR_2_0_VSS 1.71569410917e-08
R_2_14 PAR_2_0_VDD075CPU n99 0.00377712577852
C_2_14 n99 PAR_2_0_VSS 1.42757523124e-08
R_3_14 PAR_2_0_VDD075CPU n100 0.00160133993858
C_3_14 n100 PAR_2_0_VSS 6.34465159375e-08
R_4_14 PAR_2_0_VDD075CPU n101 1.47822560007
C_4_14 n101 PAR_2_0_VSS 2.82494192406e-10
R_5_14 PAR_2_0_VDD075CPU n102 3.77426174974
C_5_14 n102 PAR_2_0_VSS 2.39135912106e-10
L_6_14 PAR_2_0_VDD075CPU n103 7.36601353142e-08
R_6_14 n103 PAR_2_0_VSS 17.3275234936
G0_15 PAR_2_0_VDD075CPU PAR_0_0_VSS PAR_2_0_VDD075CPU PAR_0_0_VSS -0.599098610647
C0_15 PAR_2_0_VDD075CPU PAR_0_0_VSS 2.93630108382e-10
R_1_15 PAR_2_0_VDD075CPU n104 0.0150416980177
C_1_15 n104 PAR_0_0_VSS 9.09829198479e-10
R_2_15 PAR_2_0_VDD075CPU n105 0.304804873632
C_2_15 n105 PAR_0_0_VSS 2.55271758402e-10
L_3_15 PAR_2_0_VDD075CPU n106 4.55187229436e-10
R_3_15 n106 PAR_0_0_VSS 1.66917428573
R_4_15 PAR_2_0_VDD075CPU n107 8.79657689277
C_4_15 n107 PAR_0_0_VSS 9.07603786141e-11
R_5_15 PAR_2_0_VDD075CPU n108 43.96929905
C_5_15 n108 PAR_0_0_VSS 1.02409703002e-10
R_6_15 PAR_2_0_VDD075CPU n109 145.106882624
C_6_15 n109 PAR_0_0_VSS 1.10011264161e-10
G0_16 PAR_0_1_VSS PAR_0_0_VDD075CPU PAR_0_1_VSS PAR_0_0_VDD075CPU -0.0937306635146
C0_16 PAR_0_1_VSS PAR_0_0_VDD075CPU 1.7165145143e-10
R_1_16 PAR_0_1_VSS n110 0.0323103903056
C_1_16 n110 PAR_0_0_VDD075CPU 4.87961935102e-10
R_2_16 PAR_0_1_VSS n111 0.0311016249579
C_2_16 n111 PAR_0_0_VDD075CPU 1.65636593714e-09
R_3_16 PAR_0_1_VSS n112 0.0227681308123
C_3_16 n112 PAR_0_0_VDD075CPU 4.57247584822e-09
L_4_16 PAR_0_1_VSS n113 6.18657324247e-09
R_4_16 n113 PAR_0_0_VDD075CPU 10.6688668881
R_5_16 PAR_0_1_VSS n114 27.9957280176
C_5_16 n114 PAR_0_0_VDD075CPU 1.89239034327e-10
R_6_16 PAR_0_1_VSS n115 67.4493748962
C_6_16 n115 PAR_0_0_VDD075CPU 2.36560901271e-10
R0_17 PAR_0_1_VSS PAR_1_0_VSS 0.124606911989
C0_17 PAR_0_1_VSS PAR_1_0_VSS 1.76878829751e-10
R_1_17 PAR_0_1_VSS n116 0.414444283623
C_1_17 n116 PAR_1_0_VSS 7.62310911401e-11
R_2_17 PAR_0_1_VSS n117 0.102398436047
C_2_17 n117 PAR_1_0_VSS 2.0739939734e-09
R_3_17 PAR_0_1_VSS n118 0.414285391976
C_3_17 n118 PAR_1_0_VSS 7.60405817274e-10
R_4_17 PAR_0_1_VSS n119 0.335151229618
C_4_17 n119 PAR_1_0_VSS 2.46064973221e-09
R_5_17 PAR_0_1_VSS n120 1.54760005299
C_5_17 n120 PAR_1_0_VSS 2.69355118562e-09
R_6_17 PAR_0_1_VSS n121 3.36173913486
C_6_17 n121 PAR_1_0_VSS 4.22465927142e-09
G0_18 PAR_0_1_VSS PAR_1_0_VDD075CPU PAR_0_1_VSS PAR_1_0_VDD075CPU -0.25370974966
C0_18 PAR_0_1_VSS PAR_1_0_VDD075CPU 2.21828186408e-10
R_1_18 PAR_0_1_VSS n122 0.0892839163844
C_1_18 n122 PAR_1_0_VDD075CPU 2.80114115934e-10
R_2_18 PAR_0_1_VSS n123 0.199423100788
C_2_18 n123 PAR_1_0_VDD075CPU 3.74052338238e-10
L_3_18 PAR_0_1_VSS n124 1.65897479962e-09
R_3_18 n124 PAR_1_0_VDD075CPU 3.94151186866
R_4_18 PAR_0_1_VSS n125 23.2042390928
C_4_18 n125 PAR_1_0_VDD075CPU 3.21452468414e-10
R_5_18 PAR_0_1_VSS n126 190.690743346
C_5_18 n126 PAR_1_0_VDD075CPU 1.31663315509e-10
R0_19 PAR_0_1_VSS PAR_2_0_VSS 1468.38737402
C0_19 PAR_0_1_VSS PAR_2_0_VSS 2.36899363965e-10
R_1_19 PAR_0_1_VSS n127 0.202816417626
C_1_19 n127 PAR_2_0_VSS 1.56453371127e-10
R_2_19 PAR_0_1_VSS n128 0.665726093607
C_2_19 n128 PAR_2_0_VSS 1.56762311053e-10
R_3_19 PAR_0_1_VSS n129 0.398475158068
C_3_19 n129 PAR_2_0_VSS 6.86446828466e-10
R_4_19 PAR_0_1_VSS n130 0.179370024699
C_4_19 n130 PAR_2_0_VSS 4.68772664033e-09
R_5_19 PAR_0_1_VSS n131 1.38458894228
C_5_19 n131 PAR_2_0_VSS 3.07900660823e-09
R_6_19 PAR_0_1_VSS n132 3.01085399081
C_6_19 n132 PAR_2_0_VSS 4.74390791308e-09
G0_20 PAR_0_1_VSS PAR_2_0_VDD075CPU PAR_0_1_VSS PAR_2_0_VDD075CPU -0.1702782382
C0_20 PAR_0_1_VSS PAR_2_0_VDD075CPU 2.30582618775e-10
R_1_20 PAR_0_1_VSS n133 0.157138621904
C_1_20 n133 PAR_2_0_VDD075CPU 1.58839911535e-10
R_2_20 PAR_0_1_VSS n134 0.342575802289
C_2_20 n134 PAR_2_0_VDD075CPU 2.7109575684e-10
L_3_20 PAR_0_1_VSS n135 3.44489287708e-09
R_3_20 n135 PAR_2_0_VDD075CPU 5.87274096174
R_4_20 PAR_0_1_VSS n136 33.2522257501
C_4_20 n136 PAR_2_0_VDD075CPU 1.30797430471e-10
R_5_20 PAR_0_1_VSS n137 32.1703848881
C_5_20 n137 PAR_2_0_VDD075CPU 4.04180902142e-10
R0_21 PAR_0_1_VSS PAR_0_0_VSS 0.00414292496765
C0_21 PAR_0_1_VSS PAR_0_0_VSS 3.0152208436e-10
R_1_21 PAR_0_1_VSS n138 0.214057335734
C_1_21 n138 PAR_0_0_VSS 2.44039242493e-09
L_2_21 PAR_0_1_VSS n139 5.17070801617e-09
R_2_21 n139 PAR_0_0_VSS 0.404071767304
R0_22 PAR_0_1_VDD075CPU PAR_0_0_VDD075CPU 0.00642102539441
C0_22 PAR_0_1_VDD075CPU PAR_0_0_VDD075CPU 6.64296160007e-11
L_1_22 PAR_0_1_VDD075CPU n140 1.2820348962e-12
R_1_22 n140 PAR_0_0_VDD075CPU 0.0674276633354
L_2_22 PAR_0_1_VDD075CPU n141 3.34288418026e-12
R_2_22 n141 PAR_0_0_VDD075CPU 0.0595995388154
L_3_22 PAR_0_1_VDD075CPU n142 3.79561873444e-12
R_3_22 n142 PAR_0_0_VDD075CPU 0.0354971566435
L_4_22 PAR_0_1_VDD075CPU n143 1.38725697468e-08
R_4_22 n143 PAR_0_0_VDD075CPU 35.5453110442
L_5_22 PAR_0_1_VDD075CPU n144 2.50817085092e-07
R_5_22 n144 PAR_0_0_VDD075CPU 192.985187743
L_6_22 PAR_0_1_VDD075CPU n145 1.11753478619e-05
R_6_22 n145 PAR_0_0_VDD075CPU 1287.4939985
G0_23 PAR_0_1_VDD075CPU PAR_1_0_VSS PAR_0_1_VDD075CPU PAR_1_0_VSS -0.336222629524
C0_23 PAR_0_1_VDD075CPU PAR_1_0_VSS 1.7259942517e-10
R_1_23 PAR_0_1_VDD075CPU n146 0.28668813499
C_1_23 n146 PAR_1_0_VSS 9.87276214503e-11
R_2_23 PAR_0_1_VDD075CPU n147 0.676745121122
C_2_23 n147 PAR_1_0_VSS 1.50884102964e-10
L_3_23 PAR_0_1_VDD075CPU n148 1.20741455585e-09
R_3_23 n148 PAR_1_0_VSS 3.85378764559
L_4_23 PAR_0_1_VDD075CPU n149 2.71049708434e-08
R_4_23 n149 PAR_1_0_VSS 15.0622854471
L_5_23 PAR_0_1_VDD075CPU n150 1.06203984068e-06
R_5_23 n150 PAR_1_0_VSS 96.649477669
R0_24 PAR_0_1_VDD075CPU PAR_1_0_VDD075CPU 0.734165253428
C0_24 PAR_0_1_VDD075CPU PAR_1_0_VDD075CPU 1.69926072917e-10
L_1_24 PAR_0_1_VDD075CPU n151 5.00145631388e-12
R_1_24 n151 PAR_1_0_VDD075CPU 0.221736535841
L_2_24 PAR_0_1_VDD075CPU n152 3.53008420322e-11
R_2_24 n152 PAR_1_0_VDD075CPU 0.562638202449
L_3_24 PAR_0_1_VDD075CPU n153 3.86372017523e-10
R_3_24 n153 PAR_1_0_VDD075CPU 2.76679228653
L_4_24 PAR_0_1_VDD075CPU n154 2.40019907834e-08
R_4_24 n154 PAR_1_0_VDD075CPU 45.2589757019
L_5_24 PAR_0_1_VDD075CPU n155 1.30306918486e-06
R_5_24 n155 PAR_1_0_VDD075CPU 409.953688472
G0_25 PAR_0_1_VDD075CPU PAR_2_0_VSS PAR_0_1_VDD075CPU PAR_2_0_VSS -0.083859338916
C0_25 PAR_0_1_VDD075CPU PAR_2_0_VSS 1.92431688798e-10
R_1_25 PAR_0_1_VDD075CPU n156 3.12271630866
C_1_25 n156 PAR_2_0_VSS 3.57695977581e-11
R_2_25 PAR_0_1_VDD075CPU n157 4.3996992599
C_2_25 n157 PAR_2_0_VSS 1.12661441131e-10
L_3_25 PAR_0_1_VDD075CPU n158 2.77945914093e-08
R_3_25 n158 PAR_2_0_VSS 13.5646962706
L_4_25 PAR_0_1_VDD075CPU n159 1.19292594225e-06
R_4_25 n159 PAR_2_0_VSS 98.6333301758
G0_26 PAR_0_1_VDD075CPU PAR_2_0_VDD075CPU PAR_0_1_VDD075CPU PAR_2_0_VDD075CPU -3.57694388939
C0_26 PAR_0_1_VDD075CPU PAR_2_0_VDD075CPU 1.38157317655e-10
R_1_26 PAR_0_1_VDD075CPU n160 0.379033188374
C_1_26 n160 PAR_2_0_VDD075CPU 5.02445618041e-11
L_2_26 PAR_0_1_VDD075CPU n161 1.92652712013e-11
R_2_26 n161 PAR_2_0_VDD075CPU 0.359893827069
R_3_26 PAR_0_1_VDD075CPU n162 1.75667047938
C_3_26 n162 PAR_2_0_VDD075CPU 7.07785961104e-11
L_4_26 PAR_0_1_VDD075CPU n163 4.36978802401e-10
R_4_26 n163 PAR_2_0_VDD075CPU 1.58971743695
R_5_26 PAR_0_1_VDD075CPU n164 3.11540945015
C_5_26 n164 PAR_2_0_VDD075CPU 1.87323942936e-10
L_6_26 PAR_0_1_VDD075CPU n165 9.0042992719e-09
R_6_26 n165 PAR_2_0_VDD075CPU 6.43172541066
R_7_26 PAR_0_1_VDD075CPU n166 20.6574563941
C_7_26 n166 PAR_2_0_VDD075CPU 1.99887387758e-10
L_8_26 PAR_0_1_VDD075CPU n167 1.01920339716e-06
R_8_26 n167 PAR_2_0_VDD075CPU 71.1093706094
C0_27 PAR_0_1_VDD075CPU PAR_0_1_VSS 7.29831548902e-10
R_1_27 PAR_0_1_VDD075CPU n168 0.000954652034099
C_1_27 n168 PAR_0_1_VSS 1.78890338715e-08
R_2_27 PAR_0_1_VDD075CPU n169 0.0023371353717
C_2_27 n169 PAR_0_1_VSS 2.18829045807e-08
R_3_27 PAR_0_1_VDD075CPU n170 0.00228114412101
C_3_27 n170 PAR_0_1_VSS 4.28614223804e-08
R_4_27 PAR_0_1_VDD075CPU n171 0.504111082258
C_4_27 n171 PAR_0_1_VSS 4.11660993898e-10
R_5_27 PAR_0_1_VDD075CPU n172 27.9834545592
C_5_27 n172 PAR_0_1_VSS 5.84969571949e-11
R_6_27 PAR_0_1_VDD075CPU n173 27.5196218454
C_6_27 n173 PAR_0_1_VSS 3.33181156074e-10
G0_28 PAR_0_1_VDD075CPU PAR_0_0_VSS PAR_0_1_VDD075CPU PAR_0_0_VSS -0.847738369945
C0_28 PAR_0_1_VDD075CPU PAR_0_0_VSS 2.25651226824e-10
R_1_28 PAR_0_1_VDD075CPU n174 0.0195487494609
C_1_28 n174 PAR_0_0_VSS 7.99955770617e-10
R_2_28 PAR_0_1_VDD075CPU n175 0.122724686994
C_2_28 n175 PAR_0_0_VSS 5.48816655004e-10
R_3_28 PAR_0_1_VDD075CPU n176 0.0762112580306
C_3_28 n176 PAR_0_0_VSS 1.51454446801e-09
L_4_28 PAR_0_1_VDD075CPU n177 2.56846167091e-10
R_4_28 n177 PAR_0_0_VSS 1.17960921943
R_5_28 PAR_0_1_VDD075CPU n178 9.05621197817
C_5_28 n178 PAR_0_0_VSS 1.15536962535e-10
R_6_28 PAR_0_1_VDD075CPU n179 63.5568568794
C_6_28 n179 PAR_0_0_VSS 1.25820725423e-10
G0_29 PAR_1_1_VSS PAR_0_0_VDD075CPU PAR_1_1_VSS PAR_0_0_VDD075CPU -0.786002122851
C0_29 PAR_1_1_VSS PAR_0_0_VDD075CPU 1.19155369698e-10
L_1_29 PAR_1_1_VSS n180 3.05449766539e-11
R_1_29 n180 PAR_0_0_VDD075CPU 1.47367590068
R_2_29 PAR_1_1_VSS n181 1.41053062625
C_2_29 n181 PAR_0_0_VDD075CPU 3.35222084571e-11
R_3_29 PAR_1_1_VSS n182 24.5279510005
C_3_29 n182 PAR_0_0_VDD075CPU 5.04927461622e-12
L_4_29 PAR_1_1_VSS n183 3.70159911141e-09
R_4_29 n183 PAR_0_0_VDD075CPU 10.8760184486
R_5_29 PAR_1_1_VSS n184 29.0520415958
C_5_29 n184 PAR_0_0_VDD075CPU 2.899202419e-11
L_6_29 PAR_1_1_VSS n185 1.85871322043e-07
R_6_29 n185 PAR_0_0_VDD075CPU 64.5933996972
R_7_29 PAR_1_1_VSS n186 538.137068009
C_7_29 n186 PAR_0_0_VDD075CPU 2.42313722093e-11
R0_30 PAR_1_1_VSS PAR_1_0_VSS 0.00618777936227
C0_30 PAR_1_1_VSS PAR_1_0_VSS 4.14022732804e-11
L_1_30 PAR_1_1_VSS n187 1.6671843137e-12
R_1_30 n187 PAR_1_0_VSS 0.0752455940686
L_2_30 PAR_1_1_VSS n188 2.78635056047e-12
R_2_30 n188 PAR_1_0_VSS 0.052550276395
L_3_30 PAR_1_1_VSS n189 5.83850215663e-09
R_3_30 n189 PAR_1_0_VSS 14.8819563023
L_4_30 PAR_1_1_VSS n190 6.18336034797e-08
R_4_30 n190 PAR_1_0_VSS 29.9071854054
L_5_30 PAR_1_1_VSS n191 2.49374715404e-06
R_5_30 n191 PAR_1_0_VSS 197.21425446
G0_31 PAR_1_1_VSS PAR_1_0_VDD075CPU PAR_1_1_VSS PAR_1_0_VDD075CPU -0.065924505533
C0_31 PAR_1_1_VSS PAR_1_0_VDD075CPU 2.14160001903e-10
R_1_31 PAR_1_1_VSS n192 0.0467198009344
C_1_31 n192 PAR_1_0_VDD075CPU 3.42857223153e-10
R_2_31 PAR_1_1_VSS n193 0.0229473426528
C_2_31 n193 PAR_1_0_VDD075CPU 1.74364029994e-09
R_3_31 PAR_1_1_VSS n194 0.0524983696717
C_3_31 n194 PAR_1_0_VDD075CPU 1.14043312108e-09
L_4_31 PAR_1_1_VSS n195 3.5139158613e-09
R_4_31 n195 PAR_1_0_VDD075CPU 17.7053185721
L_5_31 PAR_1_1_VSS n196 8.37932921985e-08
R_5_31 n196 PAR_1_0_VDD075CPU 116.913917982
L_6_31 PAR_1_1_VSS n197 6.76088159711e-06
R_6_31 n197 PAR_1_0_VDD075CPU 1122.33122335
R0_32 PAR_1_1_VSS PAR_2_0_VSS 0.361033913153
C0_32 PAR_1_1_VSS PAR_2_0_VSS 1.54356248065e-10
L_1_32 PAR_1_1_VSS n198 5.09119302788e-12
R_1_32 n198 PAR_2_0_VSS 0.322933009406
L_2_32 PAR_1_1_VSS n199 2.54102011158e-11
R_2_32 n199 PAR_2_0_VSS 0.403107597387
R_3_32 PAR_1_1_VSS n200 14.2267721656
C_3_32 n200 PAR_2_0_VSS 1.27645332508e-11
R_4_32 PAR_1_1_VSS n201 7.47194914237
C_4_32 n201 PAR_2_0_VSS 7.51931782086e-11
L_5_32 PAR_1_1_VSS n202 3.94432805635e-08
R_5_32 n202 PAR_2_0_VSS 21.2943587839
L_6_32 PAR_1_1_VSS n203 1.57745090264e-06
R_6_32 n203 PAR_2_0_VSS 144.535429175
G0_33 PAR_1_1_VSS PAR_2_0_VDD075CPU PAR_1_1_VSS PAR_2_0_VDD075CPU -1.4293609722
C0_33 PAR_1_1_VSS PAR_2_0_VDD075CPU 1.28875824745e-10
L_1_33 PAR_1_1_VSS n204 1.01845470482e-11
R_1_33 n204 PAR_2_0_VDD075CPU 0.785779542036
R_2_33 PAR_1_1_VSS n205 0.793999740156
C_2_33 n205 PAR_2_0_VDD075CPU 7.6235773527e-11
R_3_33 PAR_1_1_VSS n206 8.16850502852
C_3_33 n206 PAR_2_0_VDD075CPU 1.56602712771e-11
L_4_33 PAR_1_1_VSS n207 2.30494285932e-09
R_4_33 n207 PAR_2_0_VDD075CPU 7.20753149882
R_5_33 PAR_1_1_VSS n208 21.9832096466
C_5_33 n208 PAR_2_0_VDD075CPU 3.3796221926e-11
L_6_33 PAR_1_1_VSS n209 1.51621505009e-07
R_6_33 n209 PAR_2_0_VDD075CPU 55.5690146037
R_7_33 PAR_1_1_VSS n210 498.994131028
C_7_33 n210 PAR_2_0_VDD075CPU 2.5677649857e-11
R0_34 PAR_1_1_VSS PAR_0_1_VSS 0.00382164766635
L_1_34 PAR_1_1_VSS n211 4.35996563148e-13
R_1_34 n211 PAR_0_1_VSS 0.0183636028397
L_2_34 PAR_1_1_VSS n212 2.67741251915e-12
R_2_34 n212 PAR_0_1_VSS 0.0438194591958
L_3_34 PAR_1_1_VSS n213 1.85678263293e-10
R_3_34 n213 PAR_0_1_VSS 1.30145802581
R_4_34 PAR_1_1_VSS n214 32.0067542838
C_4_34 n214 PAR_0_1_VSS 2.33623194441e-11
R_5_34 PAR_1_1_VSS n215 44.1781838327
C_5_34 n215 PAR_0_1_VSS 1.65245752358e-10
G0_35 PAR_1_1_VSS PAR_0_1_VDD075CPU PAR_1_1_VSS PAR_0_1_VDD075CPU -0.0168846490174
C0_35 PAR_1_1_VSS PAR_0_1_VDD075CPU 1.10605638454e-10
R_1_35 PAR_1_1_VSS n216 0.043675489759
C_1_35 n216 PAR_0_1_VDD075CPU 4.77200811276e-10
R_2_35 PAR_1_1_VSS n217 0.0600701467565
C_2_35 n217 PAR_0_1_VDD075CPU 8.17497407243e-10
R_3_35 PAR_1_1_VSS n218 0.222126472398
C_3_35 n218 PAR_0_1_VDD075CPU 3.61617051632e-10
L_4_35 PAR_1_1_VSS n219 2.8147934266e-08
R_4_35 n219 PAR_0_1_VDD075CPU 70.397926366
L_5_35 PAR_1_1_VSS n220 6.23490180287e-07
R_5_35 n220 PAR_0_1_VDD075CPU 442.701078445
L_6_35 PAR_1_1_VSS n221 2.29666448343e-05
R_6_35 n221 PAR_0_1_VDD075CPU 2376.27378312
R0_36 PAR_1_1_VSS PAR_0_0_VSS 0.175315789621
C0_36 PAR_1_1_VSS PAR_0_0_VSS 1.11709784576e-10
R_1_36 PAR_1_1_VSS n222 0.0184467953886
C_1_36 n222 PAR_0_0_VSS 4.71774791896e-10
L_2_36 PAR_1_1_VSS n223 2.91376870128e-11
R_2_36 n223 PAR_0_0_VSS 0.475139423028
L_3_36 PAR_1_1_VSS n224 1.08725978272e-09
R_3_36 n224 PAR_0_0_VSS 4.80264324802
R_4_36 PAR_1_1_VSS n225 14.8273350762
C_4_36 n225 PAR_0_0_VSS 7.33811465416e-11
R_5_36 PAR_1_1_VSS n226 115.903398876
C_5_36 n226 PAR_0_0_VSS 7.15935601156e-11
R0_37 PAR_1_1_VDD075CPU PAR_0_0_VDD075CPU 0.606964086843
C0_37 PAR_1_1_VDD075CPU PAR_0_0_VDD075CPU 1.3607899057e-10
L_1_37 PAR_1_1_VDD075CPU n227 5.27382455478e-12
R_1_37 n227 PAR_0_0_VDD075CPU 0.225830213092
L_2_37 PAR_1_1_VDD075CPU n228 3.43396098472e-11
R_2_37 n228 PAR_0_0_VDD075CPU 0.57038010266
L_3_37 PAR_1_1_VDD075CPU n229 6.17841823928e-10
R_3_37 n229 PAR_0_0_VDD075CPU 4.62067770062
L_4_37 PAR_1_1_VDD075CPU n230 2.56334085525e-08
R_4_37 n230 PAR_0_0_VDD075CPU 55.4838358736
L_5_37 PAR_1_1_VDD075CPU n231 6.90694291374e-07
R_5_37 n231 PAR_0_0_VDD075CPU 375.22090496
L_6_37 PAR_1_1_VDD075CPU n232 4.45253474252e-05
R_6_37 n232 PAR_0_0_VDD075CPU 2400.49039816
G0_38 PAR_1_1_VDD075CPU PAR_1_0_VSS PAR_1_1_VDD075CPU PAR_1_0_VSS -0.290781966165
C0_38 PAR_1_1_VDD075CPU PAR_1_0_VSS 1.60081945955e-10
R_1_38 PAR_1_1_VDD075CPU n233 0.106285732062
C_1_38 n233 PAR_1_0_VSS 2.25546011799e-10
R_2_38 PAR_1_1_VDD075CPU n234 0.0886367090596
C_2_38 n234 PAR_1_0_VSS 6.22745664761e-10
R_3_38 PAR_1_1_VDD075CPU n235 1.42581832124
C_3_38 n235 PAR_1_0_VSS 9.61414508437e-11
L_4_38 PAR_1_1_VDD075CPU n236 1.09948059921e-09
R_4_38 n236 PAR_1_0_VSS 4.27565466672
L_5_38 PAR_1_1_VDD075CPU n237 3.58629408953e-08
R_5_38 n237 PAR_1_0_VSS 20.5515489401
L_6_38 PAR_1_1_VDD075CPU n238 1.27412698424e-06
R_6_38 n238 PAR_1_0_VSS 121.336792068
R0_39 PAR_1_1_VDD075CPU PAR_1_0_VDD075CPU 0.00646677738992
C0_39 PAR_1_1_VDD075CPU PAR_1_0_VDD075CPU 4.33084971233e-11
L_1_39 PAR_1_1_VDD075CPU n239 9.07470864565e-13
R_1_39 n239 PAR_1_0_VDD075CPU 0.0495930356237
L_2_39 PAR_1_1_VDD075CPU n240 1.50294296351e-12
R_2_39 n240 PAR_1_0_VDD075CPU 0.0318790753645
L_3_39 PAR_1_1_VDD075CPU n241 2.58600053455e-11
R_3_39 n241 PAR_1_0_VDD075CPU 0.321833641116
L_4_39 PAR_1_1_VDD075CPU n242 6.37186245979e-09
R_4_39 n242 PAR_1_0_VDD075CPU 23.7060931565
L_5_39 PAR_1_1_VDD075CPU n243 1.23926249648e-07
R_5_39 n243 PAR_1_0_VDD075CPU 137.58868701
L_6_39 PAR_1_1_VDD075CPU n244 7.90631068507e-06
R_6_39 n244 PAR_1_0_VDD075CPU 1097.36263731
G0_40 PAR_1_1_VDD075CPU PAR_2_0_VSS PAR_1_1_VDD075CPU PAR_2_0_VSS -0.0438103406561
C0_40 PAR_1_1_VDD075CPU PAR_2_0_VSS 1.5592934328e-10
R_1_40 PAR_1_1_VDD075CPU n245 0.58622512514
C_1_40 n245 PAR_2_0_VSS 1.16309981925e-10
R_2_40 PAR_1_1_VDD075CPU n246 5.0746890019
C_2_40 n246 PAR_2_0_VSS 8.29495487991e-11
L_3_40 PAR_1_1_VDD075CPU n247 7.67773862432e-08
R_3_40 n247 PAR_2_0_VSS 22.8256600979
C0_41 PAR_1_1_VDD075CPU PAR_2_0_VDD075CPU 1.5135107399e-10
L_1_41 PAR_1_1_VDD075CPU n248 3.23295584193e-12
R_1_41 n248 PAR_2_0_VDD075CPU 0.188498893211
L_2_41 PAR_1_1_VDD075CPU n249 2.49071339255e-11
R_2_41 n249 PAR_2_0_VDD075CPU 0.418350904011
L_3_41 PAR_1_1_VDD075CPU n250 5.85040325259e-10
R_3_41 n250 PAR_2_0_VDD075CPU 4.50137529803
L_4_41 PAR_1_1_VDD075CPU n251 9.21393085377e-09
R_4_41 n251 PAR_2_0_VDD075CPU 23.3461426421
L_5_41 PAR_1_1_VDD075CPU n252 3.43628431532e-06
R_5_41 n252 PAR_2_0_VDD075CPU 2862.51273707
L_6_41 PAR_1_1_VDD075CPU n253 3.89137051059e-06
R_6_41 n253 PAR_2_0_VDD075CPU 465.399343108
G0_42 PAR_1_1_VDD075CPU PAR_0_1_VSS PAR_1_1_VDD075CPU PAR_0_1_VSS -0.0582727156659
C0_42 PAR_1_1_VDD075CPU PAR_0_1_VSS 2.25454215463e-10
R_1_42 PAR_1_1_VDD075CPU n254 0.0108659151034
C_1_42 n254 PAR_0_1_VSS 1.86754720613e-09
R_2_42 PAR_1_1_VDD075CPU n255 0.0227527342011
C_2_42 n255 PAR_0_1_VSS 2.39639198121e-09
R_3_42 PAR_1_1_VDD075CPU n256 0.204455544621
C_3_42 n256 PAR_0_1_VSS 4.77798879734e-10
L_4_42 PAR_1_1_VDD075CPU n257 8.91960086545e-09
R_4_42 n257 PAR_0_1_VSS 17.1606890916
R_5_42 PAR_1_1_VDD075CPU n258 31.4486325423
C_5_42 n258 PAR_0_1_VSS 2.4693897983e-10
R0_43 PAR_1_1_VDD075CPU PAR_0_1_VDD075CPU 0.00449240814966
C0_43 PAR_1_1_VDD075CPU PAR_0_1_VDD075CPU 2.85602435421e-12
L_1_43 PAR_1_1_VDD075CPU n259 3.61602711007e-13
R_1_43 n259 PAR_0_1_VDD075CPU 0.01848730864
L_2_43 PAR_1_1_VDD075CPU n260 1.69479194567e-12
R_2_43 n260 PAR_0_1_VDD075CPU 0.033508808423
L_3_43 PAR_1_1_VDD075CPU n261 1.56405548166e-11
R_3_43 n261 PAR_0_1_VDD075CPU 0.175917094732
L_4_43 PAR_1_1_VDD075CPU n262 9.03004024225e-09
R_4_43 n262 PAR_0_1_VDD075CPU 29.8493814516
L_5_43 PAR_1_1_VDD075CPU n263 3.12086185914e-07
R_5_43 n263 PAR_0_1_VDD075CPU 238.900756672
L_6_43 PAR_1_1_VDD075CPU n264 9.47309075963e-05
R_6_43 n264 PAR_0_1_VDD075CPU 4639.76068302
G0_44 PAR_1_1_VDD075CPU PAR_1_1_VSS PAR_1_1_VDD075CPU PAR_1_1_VSS -0.0074657374646
C0_44 PAR_1_1_VDD075CPU PAR_1_1_VSS 3.44432247418e-10
R_1_44 PAR_1_1_VDD075CPU n265 0.000880678038436
C_1_44 n265 PAR_1_1_VSS 1.32061354983e-08
R_2_44 PAR_1_1_VDD075CPU n266 0.0018960547037
C_2_44 n266 PAR_1_1_VSS 1.5826372757e-08
R_3_44 PAR_1_1_VDD075CPU n267 0.00358563369228
C_3_44 n267 PAR_1_1_VSS 1.55618609428e-08
R_4_44 PAR_1_1_VDD075CPU n268 0.0116393794218
C_4_44 n268 PAR_1_1_VSS 8.02068820895e-09
L_5_44 PAR_1_1_VDD075CPU n269 9.06542071097e-08
R_5_44 n269 PAR_1_1_VSS 147.617454155
L_6_44 PAR_1_1_VDD075CPU n270 7.14348497621e-06
R_6_44 n270 PAR_1_1_VSS 1446.18797926
G0_45 PAR_1_1_VDD075CPU PAR_0_0_VSS PAR_1_1_VDD075CPU PAR_0_0_VSS -0.215624106389
C0_45 PAR_1_1_VDD075CPU PAR_0_0_VSS 1.87079167157e-10
R_1_45 PAR_1_1_VDD075CPU n271 0.0240156688224
C_1_45 n271 PAR_0_0_VSS 5.17926096787e-10
R_2_45 PAR_1_1_VDD075CPU n272 0.882098664494
C_2_45 n272 PAR_0_0_VSS 6.67102133527e-11
L_3_45 PAR_1_1_VDD075CPU n273 1.2851246403e-09
R_3_45 n273 PAR_0_0_VSS 4.63770032368
R_4_45 PAR_1_1_VDD075CPU n274 10.6773476741
C_4_45 n274 PAR_0_0_VSS 8.72676685053e-11
R_5_45 PAR_1_1_VDD075CPU n275 86.9268275311
C_5_45 n275 PAR_0_0_VSS 5.09522180945e-11
R_6_45 PAR_1_1_VDD075CPU n276 265.676756268
C_6_45 n276 PAR_0_0_VSS 5.80736670196e-11
G0_46 PAR_2_1_VSS PAR_0_0_VDD075CPU PAR_2_1_VSS PAR_0_0_VDD075CPU -1.57334440423
C0_46 PAR_2_1_VSS PAR_0_0_VDD075CPU 1.33221135017e-10
R_1_46 PAR_2_1_VSS n277 2.03581420002
C_1_46 n277 PAR_0_0_VDD075CPU 1.3297666991e-11
L_2_46 PAR_2_1_VSS n278 1.07459968232e-10
R_2_46 n278 PAR_0_0_VDD075CPU 0.807186547584
R_3_46 PAR_2_1_VSS n279 1.01137909461
C_3_46 n279 PAR_0_0_VDD075CPU 2.06891618559e-10
L_4_46 PAR_2_1_VSS n280 2.46557284128e-09
R_4_46 n280 PAR_0_0_VDD075CPU 3.37319505794
R_5_46 PAR_2_1_VSS n281 10.7076113915
C_5_46 n281 PAR_0_0_VDD075CPU 2.50018853197e-10
L_6_46 PAR_2_1_VSS n282 3.23064472369e-07
R_6_46 n282 PAR_0_0_VDD075CPU 26.3029330659
R0_47 PAR_2_1_VSS PAR_1_0_VSS 0.17907171236
C0_47 PAR_2_1_VSS PAR_1_0_VSS 1.64961727667e-10
R_1_47 PAR_2_1_VSS n283 0.473714602388
C_1_47 n283 PAR_1_0_VSS 3.58086703367e-11
L_2_47 PAR_2_1_VSS n284 3.61807140524e-11
R_2_47 n284 PAR_1_0_VSS 0.515161440967
R_3_47 PAR_2_1_VSS n285 0.435603020982
C_3_47 n285 PAR_1_0_VSS 5.07631617533e-10
R_4_47 PAR_2_1_VSS n286 1.11151322175
C_4_47 n286 PAR_1_0_VSS 6.72169132872e-10
L_5_47 PAR_2_1_VSS n287 3.00576262324e-08
R_5_47 n287 PAR_1_0_VSS 8.36268774098
L_6_47 PAR_2_1_VSS n288 3.1221078081e-07
R_6_47 n288 PAR_1_0_VSS 22.9816077475
G0_48 PAR_2_1_VSS PAR_1_0_VDD075CPU PAR_2_1_VSS PAR_1_0_VDD075CPU -0.111143516258
C0_48 PAR_2_1_VSS PAR_1_0_VDD075CPU 1.83547661967e-10
R_1_48 PAR_2_1_VSS n289 0.230067374025
C_1_48 n289 PAR_1_0_VDD075CPU 2.28989943062e-10
R_2_48 PAR_2_1_VSS n290 0.854714965837
C_2_48 n290 PAR_1_0_VDD075CPU 9.73687496416e-11
L_3_48 PAR_2_1_VSS n291 3.43066928765e-09
R_3_48 n291 PAR_1_0_VDD075CPU 13.3424401936
L_4_48 PAR_2_1_VSS n292 3.31724344138e-08
R_4_48 n292 PAR_1_0_VDD075CPU 40.4328966428
L_5_48 PAR_2_1_VSS n293 3.981882961e-07
R_5_48 n293 PAR_1_0_VDD075CPU 122.447356404
L_6_48 PAR_2_1_VSS n294 3.96359196668e-06
R_6_48 n294 PAR_1_0_VDD075CPU 303.435008761
R0_49 PAR_2_1_VSS PAR_2_0_VSS 0.00633883681869
C0_49 PAR_2_1_VSS PAR_2_0_VSS 1.25444406711e-10
L_1_49 PAR_2_1_VSS n295 4.676058016e-13
R_1_49 n295 PAR_2_0_VSS 0.0237350772655
L_2_49 PAR_2_1_VSS n296 4.8056210426e-12
R_2_49 n296 PAR_2_0_VSS 0.0467083904877
R_3_49 PAR_2_1_VSS n297 0.602751333083
C_3_49 n297 PAR_2_0_VSS 1.22332971895e-09
L_4_49 PAR_2_1_VSS n298 4.28961975198e-08
R_4_49 n298 PAR_2_0_VSS 6.65613608616
G0_50 PAR_2_1_VSS PAR_2_0_VDD075CPU PAR_2_1_VSS PAR_2_0_VDD075CPU -0.0576523244936
C0_50 PAR_2_1_VSS PAR_2_0_VDD075CPU 1.49510256948e-10
R_1_50 PAR_2_1_VSS n299 0.0115508429002
C_1_50 n299 PAR_2_0_VDD075CPU 1.41026462201e-09
R_2_50 PAR_2_1_VSS n300 0.0974951901073
C_2_50 n300 PAR_2_0_VDD075CPU 5.19486285377e-10
R_3_50 PAR_2_1_VSS n301 0.0255180120061
C_3_50 n301 PAR_2_0_VDD075CPU 4.09317585767e-09
L_4_50 PAR_2_1_VSS n302 1.63922907148e-08
R_4_50 n302 PAR_2_0_VDD075CPU 25.1300454164
L_5_50 PAR_2_1_VSS n303 1.82226778978e-07
R_5_50 n303 PAR_2_0_VDD075CPU 77.7507155254
L_6_50 PAR_2_1_VSS n304 2.25968497396e-06
R_6_50 n304 PAR_2_0_VDD075CPU 200.091843439
R0_51 PAR_2_1_VSS PAR_0_1_VSS 126603.284989
C0_51 PAR_2_1_VSS PAR_0_1_VSS 1.74841548134e-10
R_1_51 PAR_2_1_VSS n305 0.247254728459
C_1_51 n305 PAR_0_1_VSS 1.08643412883e-10
R_2_51 PAR_2_1_VSS n306 0.557364750136
C_2_51 n306 PAR_0_1_VSS 3.4241212634e-10
R_3_51 PAR_2_1_VSS n307 0.790131064169
C_3_51 n307 PAR_0_1_VSS 4.88601988956e-10
R_4_51 PAR_2_1_VSS n308 2.13223877735
C_4_51 n308 PAR_0_1_VSS 4.66200487282e-10
R_5_51 PAR_2_1_VSS n309 3.38133902923
C_5_51 n309 PAR_0_1_VSS 1.14474597793e-09
R_6_51 PAR_2_1_VSS n310 9.02969107983
C_6_51 n310 PAR_0_1_VSS 1.54482794269e-09
G0_52 PAR_2_1_VSS PAR_0_1_VDD075CPU PAR_2_1_VSS PAR_0_1_VDD075CPU -2.74032878782
C0_52 PAR_2_1_VSS PAR_0_1_VDD075CPU 1.14880458296e-10
R_1_52 PAR_2_1_VSS n311 1.06680957336
C_1_52 n311 PAR_0_1_VDD075CPU 1.82472500137e-11
L_2_52 PAR_2_1_VSS n312 3.10891653121e-11
R_2_52 n312 PAR_0_1_VDD075CPU 0.459599630207
R_3_52 PAR_2_1_VSS n313 0.603933739823
C_3_52 n313 PAR_0_1_VDD075CPU 1.75895108712e-10
L_4_52 PAR_2_1_VSS n314 4.52602306406e-10
R_4_52 n314 PAR_0_1_VDD075CPU 2.11722140213
R_5_52 PAR_2_1_VSS n315 8.00803807784
C_5_52 n315 PAR_0_1_VDD075CPU 7.15150731428e-11
L_6_52 PAR_2_1_VSS n316 1.74457507881e-08
R_6_52 n316 PAR_0_1_VDD075CPU 12.1239751059
R_7_52 PAR_2_1_VSS n317 44.9053606746
C_7_52 n317 PAR_0_1_VDD075CPU 9.17937160748e-11
L_8_52 PAR_2_1_VSS n318 1.46027081675e-06
R_8_52 n318 PAR_0_1_VDD075CPU 102.842219808
R0_53 PAR_2_1_VSS PAR_1_1_VSS 0.00485917844921
C0_53 PAR_2_1_VSS PAR_1_1_VSS 2.38267679943e-11
L_1_53 PAR_2_1_VSS n319 2.54039145528e-13
R_1_53 n319 PAR_1_1_VSS 0.0125186676337
L_2_53 PAR_2_1_VSS n320 2.19681157585e-12
R_2_53 n320 PAR_1_1_VSS 0.040416824622
L_3_53 PAR_2_1_VSS n321 8.27708525021e-12
R_3_53 n321 PAR_1_1_VSS 0.08503521595
L_4_53 PAR_2_1_VSS n322 2.28427260441e-08
R_4_53 n322 PAR_1_1_VSS 53.8831750137
L_5_53 PAR_2_1_VSS n323 2.39014623564e-07
R_5_53 n323 PAR_1_1_VSS 139.767613704
L_6_53 PAR_2_1_VSS n324 3.57187373453e-06
R_6_53 n324 PAR_1_1_VSS 374.45570166
G0_54 PAR_2_1_VSS PAR_1_1_VDD075CPU PAR_2_1_VSS PAR_1_1_VDD075CPU -0.0191266237518
C0_54 PAR_2_1_VSS PAR_1_1_VDD075CPU 1.12950961305e-10
R_1_54 PAR_2_1_VSS n325 0.00781956803086
C_1_54 n325 PAR_1_1_VDD075CPU 2.45599867972e-09
R_2_54 PAR_2_1_VSS n326 0.0302800069405
C_2_54 n326 PAR_1_1_VDD075CPU 1.7457468222e-09
R_3_54 PAR_2_1_VSS n327 0.0659577420819
C_3_54 n327 PAR_1_1_VDD075CPU 1.43793027525e-09
L_4_54 PAR_2_1_VSS n328 6.1804153016e-08
R_4_54 n328 PAR_1_1_VDD075CPU 83.6630299251
L_5_54 PAR_2_1_VSS n329 6.19946092957e-07
R_5_54 n329 PAR_1_1_VDD075CPU 195.227099046
L_6_54 PAR_2_1_VSS n330 6.29142542693e-06
R_6_54 n330 PAR_1_1_VDD075CPU 487.40646702
R0_55 PAR_2_1_VSS PAR_0_0_VSS 542938.032846
C0_55 PAR_2_1_VSS PAR_0_0_VSS 2.49503397437e-10
R_1_55 PAR_2_1_VSS n331 0.0244924388719
C_1_55 n331 PAR_0_0_VSS 6.23467044988e-10
R_2_55 PAR_2_1_VSS n332 0.276443081583
C_2_55 n332 PAR_0_0_VSS 6.61201906815e-10
R_3_55 PAR_2_1_VSS n333 0.622255421563
C_3_55 n333 PAR_0_0_VSS 5.97288231886e-10
R_4_55 PAR_2_1_VSS n334 0.526829921341
C_4_55 n334 PAR_0_0_VSS 2.03797680075e-09
R_5_55 PAR_2_1_VSS n335 1.78661692727
C_5_55 n335 PAR_0_0_VSS 1.4742744145e-09
R_6_55 PAR_2_1_VSS n336 21.7985908427
C_6_55 n336 PAR_0_0_VSS 5.86980225826e-10
G0_56 PAR_2_1_VDD075CPU PAR_0_0_VDD075CPU PAR_2_1_VDD075CPU PAR_0_0_VDD075CPU -1.50862676482
C0_56 PAR_2_1_VDD075CPU PAR_0_0_VDD075CPU 1.00094719388e-10
R_1_56 PAR_2_1_VDD075CPU n337 0.918602417685
C_1_56 n337 PAR_0_0_VDD075CPU 2.64894997594e-11
L_2_56 PAR_2_1_VDD075CPU n338 9.71819426107e-11
R_2_56 n338 PAR_0_0_VDD075CPU 0.779698549632
R_3_56 PAR_2_1_VDD075CPU n339 2.54967574448
C_3_56 n339 PAR_0_0_VDD075CPU 1.7041228404e-10
L_4_56 PAR_2_1_VDD075CPU n340 6.15998346647e-09
R_4_56 n340 PAR_0_0_VDD075CPU 4.42328025522
R_5_56 PAR_2_1_VDD075CPU n341 35.9585629145
C_5_56 n341 PAR_0_0_VDD075CPU 2.48381685309e-10
G0_57 PAR_2_1_VDD075CPU PAR_1_0_VSS PAR_2_1_VDD075CPU PAR_1_0_VSS -0.434624701574
C0_57 PAR_2_1_VDD075CPU PAR_1_0_VSS 1.62164065416e-10
R_1_57 PAR_2_1_VDD075CPU n342 0.353258267855
C_1_57 n342 PAR_1_0_VSS 7.99306767763e-11
R_2_57 PAR_2_1_VDD075CPU n343 0.461326778037
C_2_57 n343 PAR_1_0_VSS 2.14050852978e-10
L_3_57 PAR_2_1_VDD075CPU n344 8.44833089065e-10
R_3_57 n344 PAR_1_0_VSS 2.82371103721
L_4_57 PAR_2_1_VDD075CPU n345 2.36289339548e-08
R_4_57 n345 PAR_1_0_VSS 14.2327218157
L_5_57 PAR_2_1_VDD075CPU n346 1.02434750024e-06
R_5_57 n346 PAR_1_0_VSS 97.8455585959
R0_58 PAR_2_1_VDD075CPU PAR_1_0_VDD075CPU 1.15706428935
C0_58 PAR_2_1_VDD075CPU PAR_1_0_VDD075CPU 1.62016949441e-10
L_1_58 PAR_2_1_VDD075CPU n347 4.24364907862e-12
R_1_58 n347 PAR_1_0_VDD075CPU 0.210491545946
L_2_58 PAR_2_1_VDD075CPU n348 3.2891087828e-11
R_2_58 n348 PAR_1_0_VDD075CPU 0.530433132776
L_3_58 PAR_2_1_VDD075CPU n349 2.5929945852e-10
R_3_58 n349 PAR_1_0_VDD075CPU 1.96109064702
L_4_58 PAR_2_1_VDD075CPU n350 2.33541006039e-08
R_4_58 n350 PAR_1_0_VDD075CPU 46.603170444
L_5_58 PAR_2_1_VDD075CPU n351 8.72852553529e-07
R_5_58 n351 PAR_1_0_VDD075CPU 373.752307606
L_6_58 PAR_2_1_VDD075CPU n352 6.58919320108e-05
R_6_58 n352 PAR_1_0_VDD075CPU 2289.69278334
G0_59 PAR_2_1_VDD075CPU PAR_2_0_VSS PAR_2_1_VDD075CPU PAR_2_0_VSS -0.102798376386
C0_59 PAR_2_1_VDD075CPU PAR_2_0_VSS 1.54888138013e-10
R_1_59 PAR_2_1_VDD075CPU n353 0.0511041302243
C_1_59 n353 PAR_2_0_VSS 4.31004347541e-10
R_2_59 PAR_2_1_VDD075CPU n354 0.674634918727
C_2_59 n354 PAR_2_0_VSS 1.01365226278e-10
R_3_59 PAR_2_1_VDD075CPU n355 0.0718352577989
C_3_59 n355 PAR_2_0_VSS 1.52915010504e-09
R_4_59 PAR_2_1_VDD075CPU n356 5.21335047362
C_4_59 n356 PAR_2_0_VSS 1.08133968727e-10
L_5_59 PAR_2_1_VDD075CPU n357 1.84294799193e-08
R_5_59 n357 PAR_2_0_VSS 10.9625281566
L_6_59 PAR_2_1_VDD075CPU n358 8.97520957947e-07
R_6_59 n358 PAR_2_0_VSS 86.3666394317
R0_60 PAR_2_1_VDD075CPU PAR_2_0_VDD075CPU 0.00743106565858
C0_60 PAR_2_1_VDD075CPU PAR_2_0_VDD075CPU 1.15402665617e-10
L_1_60 PAR_2_1_VDD075CPU n359 3.51044871528e-13
R_1_60 n359 PAR_2_0_VDD075CPU 0.0193009506274
L_2_60 PAR_2_1_VDD075CPU n360 9.79627871611e-12
R_2_60 n360 PAR_2_0_VDD075CPU 0.178162270406
L_3_60 PAR_2_1_VDD075CPU n361 3.86906992649e-12
R_3_60 n361 PAR_2_0_VDD075CPU 0.0361217455753
L_4_60 PAR_2_1_VDD075CPU n362 8.152471535e-09
R_4_60 n362 PAR_2_0_VDD075CPU 22.7205720064
L_5_60 PAR_2_1_VDD075CPU n363 1.45389943285e-07
R_5_60 n363 PAR_2_0_VDD075CPU 133.685546421
L_6_60 PAR_2_1_VDD075CPU n364 7.13276458253e-06
R_6_60 n364 PAR_2_0_VDD075CPU 910.431598717
G0_61 PAR_2_1_VDD075CPU PAR_0_1_VSS PAR_2_1_VDD075CPU PAR_0_1_VSS -0.235083426456
C0_61 PAR_2_1_VDD075CPU PAR_0_1_VSS 1.52926795705e-10
R_1_61 PAR_2_1_VDD075CPU n365 0.202023805349
C_1_61 n365 PAR_0_1_VSS 9.99689205674e-11
R_2_61 PAR_2_1_VDD075CPU n366 0.408270094669
C_2_61 n366 PAR_0_1_VSS 2.15500620609e-10
L_3_61 PAR_2_1_VDD075CPU n367 1.67935697479e-09
R_3_61 n367 PAR_0_1_VSS 4.25380897286
R_4_61 PAR_2_1_VDD075CPU n368 29.2976113465
C_4_61 n368 PAR_0_1_VSS 3.04190907029e-10
G0_62 PAR_2_1_VDD075CPU PAR_0_1_VDD075CPU PAR_2_1_VDD075CPU PAR_0_1_VDD075CPU -2.00552979228
C0_62 PAR_2_1_VDD075CPU PAR_0_1_VDD075CPU 9.49496702295e-11
R_1_62 PAR_2_1_VDD075CPU n369 0.526877342246
C_1_62 n369 PAR_0_1_VDD075CPU 3.69564924576e-11
L_2_62 PAR_2_1_VDD075CPU n370 2.75521662017e-11
R_2_62 n370 PAR_0_1_VDD075CPU 0.561069091901
R_3_62 PAR_2_1_VDD075CPU n371 49.1817445374
C_3_62 n371 PAR_0_1_VDD075CPU 2.60200710284e-12
L_4_62 PAR_2_1_VDD075CPU n372 1.89612624616e-09
R_4_62 n372 PAR_0_1_VDD075CPU 5.32514359365
R_5_62 PAR_2_1_VDD075CPU n373 12.1620422601
C_5_62 n373 PAR_0_1_VDD075CPU 7.30506494313e-11
L_6_62 PAR_2_1_VDD075CPU n374 8.46625066742e-08
R_6_62 n374 PAR_0_1_VDD075CPU 28.3934490008
R_7_62 PAR_2_1_VDD075CPU n375 200.037738994
C_7_62 n375 PAR_0_1_VDD075CPU 6.56692465283e-11
G0_63 PAR_2_1_VDD075CPU PAR_1_1_VSS PAR_2_1_VDD075CPU PAR_1_1_VSS -0.0183018553785
C0_63 PAR_2_1_VDD075CPU PAR_1_1_VSS 7.20515548552e-11
R_1_63 PAR_2_1_VDD075CPU n376 0.0238110361167
C_1_63 n376 PAR_1_1_VSS 9.78020024667e-10
R_2_63 PAR_2_1_VDD075CPU n377 0.0904025228076
C_2_63 n377 PAR_1_1_VSS 6.39274326846e-10
R_3_63 PAR_2_1_VDD075CPU n378 0.164496358824
C_3_63 n378 PAR_1_1_VSS 5.8941466328e-10
L_4_63 PAR_2_1_VDD075CPU n379 2.30004058165e-08
R_4_63 n379 PAR_1_1_VSS 65.7306164894
L_5_63 PAR_2_1_VDD075CPU n380 4.24433511997e-07
R_5_63 n380 PAR_1_1_VSS 379.215417902
L_6_63 PAR_2_1_VDD075CPU n381 1.90288749065e-05
R_6_63 n381 PAR_1_1_VSS 2216.19633142
R0_64 PAR_2_1_VDD075CPU PAR_1_1_VDD075CPU 0.00519092338245
C0_64 PAR_2_1_VDD075CPU PAR_1_1_VDD075CPU 4.30806693832e-11
L_1_64 PAR_2_1_VDD075CPU n382 2.43602498945e-13
R_1_64 n382 PAR_1_1_VDD075CPU 0.0118342551808
L_2_64 PAR_2_1_VDD075CPU n383 3.07750439338e-12
R_2_64 n383 PAR_1_1_VDD075CPU 0.0553309149764
L_3_64 PAR_2_1_VDD075CPU n384 1.24964618136e-11
R_3_64 n384 PAR_1_1_VDD075CPU 0.128133545175
L_4_64 PAR_2_1_VDD075CPU n385 1.49672524823e-08
R_4_64 n385 PAR_1_1_VDD075CPU 42.2722803563
L_5_64 PAR_2_1_VDD075CPU n386 4.04751462451e-07
R_5_64 n386 PAR_1_1_VDD075CPU 273.341487283
L_6_64 PAR_2_1_VDD075CPU n387 5.41988279437e-05
R_6_64 n387 PAR_1_1_VDD075CPU 2490.32189585
G0_65 PAR_2_1_VDD075CPU PAR_2_1_VSS PAR_2_1_VDD075CPU PAR_2_1_VSS -0.00164315312782
C0_65 PAR_2_1_VDD075CPU PAR_2_1_VSS 2.98762207882e-10
R_1_65 PAR_2_1_VDD075CPU n388 0.000696467104255
C_1_65 n388 PAR_2_1_VSS 2.35769089626e-08
R_2_65 PAR_2_1_VDD075CPU n389 0.00475334903745
C_2_65 n389 PAR_2_1_VSS 1.08661891386e-08
R_3_65 PAR_2_1_VDD075CPU n390 0.00262156431552
C_3_65 n390 PAR_2_1_VSS 3.88523932418e-08
R_4_65 PAR_2_1_VDD075CPU n391 0.440029435983
C_4_65 n391 PAR_2_1_VSS 5.26509723306e-10
R_5_65 PAR_2_1_VDD075CPU n392 2.37180696753
C_5_65 n392 PAR_2_1_VSS 6.21100123963e-10
L_6_65 PAR_2_1_VDD075CPU n393 1.31238791419e-05
R_6_65 n393 PAR_2_1_VSS 608.585080421
G0_66 PAR_2_1_VDD075CPU PAR_0_0_VSS PAR_2_1_VDD075CPU PAR_0_0_VSS -0.859048054364
C0_66 PAR_2_1_VDD075CPU PAR_0_0_VSS 1.87761779357e-10
R_1_66 PAR_2_1_VDD075CPU n394 0.0204765233455
C_1_66 n394 PAR_0_0_VSS 6.34461229823e-10
R_2_66 PAR_2_1_VDD075CPU n395 0.342764009115
C_2_66 n395 PAR_0_0_VSS 2.37009334331e-10
L_3_66 PAR_2_1_VDD075CPU n396 2.79004137791e-10
R_3_66 n396 PAR_0_0_VSS 1.16407922913
R_4_66 PAR_2_1_VDD075CPU n397 15.6011181698
C_4_66 n397 PAR_0_0_VSS 6.73721065156e-11
R_5_66 PAR_2_1_VDD075CPU n398 86.33335089
C_5_66 n398 PAR_0_0_VSS 1.07027704277e-10
G0_67 PAR_0_2_VSS PAR_0_0_VDD075CPU PAR_0_2_VSS PAR_0_0_VDD075CPU -0.356424303917
C0_67 PAR_0_2_VSS PAR_0_0_VDD075CPU 1.77783459581e-10
R_1_67 PAR_0_2_VSS n399 0.117452719302
C_1_67 n399 PAR_0_0_VDD075CPU 1.49693625377e-10
R_2_67 PAR_0_2_VSS n400 0.366350906281
C_2_67 n400 PAR_0_0_VDD075CPU 2.16405302777e-10
L_3_67 PAR_0_2_VSS n401 8.58800450478e-10
R_3_67 n401 PAR_0_0_VDD075CPU 3.44213908233
L_4_67 PAR_0_2_VSS n402 1.19718590284e-08
R_4_67 n402 PAR_0_0_VDD075CPU 15.1728299052
R_5_67 PAR_0_2_VSS n403 29.8178439809
C_5_67 n403 PAR_0_0_VDD075CPU 1.74548809288e-10
R_6_67 PAR_0_2_VSS n404 69.6808467889
C_6_67 n404 PAR_0_0_VDD075CPU 2.19780597827e-10
R0_68 PAR_0_2_VSS PAR_1_0_VSS 60.3559741841
C0_68 PAR_0_2_VSS PAR_1_0_VSS 1.76457499001e-10
R_1_68 PAR_0_2_VSS n405 0.284205275965
C_1_68 n405 PAR_1_0_VSS 1.2181132164e-10
R_2_68 PAR_0_2_VSS n406 0.3478970299
C_2_68 n406 PAR_1_0_VSS 4.40811216739e-10
R_3_68 PAR_0_2_VSS n407 0.120102046524
C_3_68 n407 PAR_1_0_VSS 2.01726837851e-09
R_4_68 PAR_0_2_VSS n408 0.320162303304
C_4_68 n408 PAR_1_0_VSS 2.52224638204e-09
R_5_68 PAR_0_2_VSS n409 1.5305476949
C_5_68 n409 PAR_1_0_VSS 2.94359200102e-09
R_6_68 PAR_0_2_VSS n410 3.61995766301
C_6_68 n410 PAR_1_0_VSS 3.94652590357e-09
G0_69 PAR_0_2_VSS PAR_1_0_VDD075CPU PAR_0_2_VSS PAR_1_0_VDD075CPU -0.267838927872
C0_69 PAR_0_2_VSS PAR_1_0_VDD075CPU 2.00193726743e-10
R_1_69 PAR_0_2_VSS n411 0.188642782805
C_1_69 n411 PAR_1_0_VDD075CPU 1.13865828951e-10
R_2_69 PAR_0_2_VSS n412 0.343225422593
C_2_69 n412 PAR_1_0_VDD075CPU 2.33616951353e-10
L_3_69 PAR_0_2_VSS n413 1.34700675259e-09
R_3_69 n413 PAR_1_0_VDD075CPU 4.07933139289
L_4_69 PAR_0_2_VSS n414 7.00484023577e-08
R_4_69 n414 PAR_1_0_VDD075CPU 44.0514669019
R_5_69 PAR_0_2_VSS n415 18.189792175
C_5_69 n415 PAR_1_0_VDD075CPU 3.94576724616e-10
R0_70 PAR_0_2_VSS PAR_2_0_VSS 3490.09148369
C0_70 PAR_0_2_VSS PAR_2_0_VSS 2.22691160557e-10
R_1_70 PAR_0_2_VSS n416 0.23456727038
C_1_70 n416 PAR_2_0_VSS 1.30749120901e-10
R_2_70 PAR_0_2_VSS n417 0.605001105193
C_2_70 n417 PAR_2_0_VSS 1.58934016311e-10
R_3_70 PAR_0_2_VSS n418 0.463281668475
C_3_70 n418 PAR_2_0_VSS 5.50997055297e-10
R_4_70 PAR_0_2_VSS n419 0.188561672577
C_4_70 n419 PAR_2_0_VSS 4.53847580328e-09
R_5_70 PAR_0_2_VSS n420 1.42679892091
C_5_70 n420 PAR_2_0_VSS 3.29324892717e-09
R_6_70 PAR_0_2_VSS n421 3.51428755351
C_6_70 n421 PAR_2_0_VSS 4.13829638545e-09
G0_71 PAR_0_2_VSS PAR_2_0_VDD075CPU PAR_0_2_VSS PAR_2_0_VDD075CPU -0.12116343972
C0_71 PAR_0_2_VSS PAR_2_0_VDD075CPU 2.14097884515e-10
R_1_71 PAR_0_2_VSS n422 0.172082931645
C_1_71 n422 PAR_2_0_VDD075CPU 1.35506356322e-10
R_2_71 PAR_0_2_VSS n423 0.343049109844
C_2_71 n423 PAR_2_0_VDD075CPU 2.51890758125e-10
L_3_71 PAR_0_2_VSS n424 5.1296349708e-09
R_3_71 n424 PAR_2_0_VDD075CPU 8.25331452265
R_4_71 PAR_0_2_VSS n425 21.7724297109
C_4_71 n425 PAR_2_0_VDD075CPU 2.78844961842e-10
R_5_71 PAR_0_2_VSS n426 74.669581611
C_5_71 n426 PAR_2_0_VDD075CPU 2.30114817779e-10
R0_72 PAR_0_2_VSS PAR_0_1_VSS 0.00481653905856
L_1_72 PAR_0_2_VSS n427 4.68527487456e-12
R_1_72 n427 PAR_0_1_VSS 0.0489619243562
L_2_72 PAR_0_2_VSS n428 2.31755618691e-10
R_2_72 n428 PAR_0_1_VSS 0.245339245001
L_3_72 PAR_0_2_VSS n429 1.18175208038e-09
R_3_72 n429 PAR_0_1_VSS 0.30738415642
L_4_72 PAR_0_2_VSS n430 2.52120717145e-08
R_4_72 n430 PAR_0_1_VSS 2.01906378175
G0_73 PAR_0_2_VSS PAR_0_1_VDD075CPU PAR_0_2_VSS PAR_0_1_VDD075CPU -0.0566736518668
C0_73 PAR_0_2_VSS PAR_0_1_VDD075CPU 1.56314094473e-10
R_1_73 PAR_0_2_VSS n431 0.135485450751
C_1_73 n431 PAR_0_1_VDD075CPU 1.70046202555e-10
R_2_73 PAR_0_2_VSS n432 0.0586665919115
C_2_73 n432 PAR_0_1_VDD075CPU 1.80753293857e-09
L_3_73 PAR_0_2_VSS n433 6.83511945502e-09
R_3_73 n433 PAR_0_1_VDD075CPU 17.6448828957
R_4_73 PAR_0_2_VSS n434 28.6306974444
C_4_73 n434 PAR_0_1_VDD075CPU 1.89861283111e-10
R_5_73 PAR_0_2_VSS n435 91.4460146561
C_5_73 n435 PAR_0_1_VDD075CPU 1.79165555381e-10
R0_74 PAR_0_2_VSS PAR_1_1_VSS 0.141678167332
C0_74 PAR_0_2_VSS PAR_1_1_VSS 1.19732124955e-10
R_1_74 PAR_0_2_VSS n436 0.447569126139
C_1_74 n436 PAR_1_1_VSS 4.46036375659e-11
R_2_74 PAR_0_2_VSS n437 1.29936927092
C_2_74 n437 PAR_1_1_VSS 4.11652212476e-11
L_3_74 PAR_0_2_VSS n438 1.06614229381e-10
R_3_74 n438 PAR_1_1_VSS 0.997957118749
L_4_74 PAR_0_2_VSS n439 2.87454766895e-08
R_4_74 n439 PAR_1_1_VSS 44.0156562085
R_5_74 PAR_0_2_VSS n440 51.8588154557
C_5_74 n440 PAR_1_1_VSS 9.95079831306e-11
R_6_74 PAR_0_2_VSS n441 133.91962976
C_6_74 n441 PAR_1_1_VSS 1.16592759349e-10
G0_75 PAR_0_2_VSS PAR_1_1_VDD075CPU PAR_0_2_VSS PAR_1_1_VDD075CPU -0.0307514315381
C0_75 PAR_0_2_VSS PAR_1_1_VDD075CPU 1.3648021945e-10
R_1_75 PAR_0_2_VSS n442 0.344231606017
C_1_75 n442 PAR_1_1_VDD075CPU 7.60877962218e-11
R_2_75 PAR_0_2_VSS n443 0.464192816726
C_2_75 n443 PAR_1_1_VDD075CPU 2.1303065537e-10
L_3_75 PAR_0_2_VSS n444 2.16904367927e-08
R_3_75 n444 PAR_1_1_VDD075CPU 32.5188084423
R_4_75 PAR_0_2_VSS n445 41.0286210767
C_4_75 n445 PAR_1_1_VDD075CPU 1.26356199592e-10
R_5_75 PAR_0_2_VSS n446 108.449293138
C_5_75 n446 PAR_1_1_VDD075CPU 1.45342439766e-10
R0_76 PAR_0_2_VSS PAR_2_1_VSS 68506.692799
C0_76 PAR_0_2_VSS PAR_2_1_VSS 1.65868630785e-10
R_1_76 PAR_0_2_VSS n447 0.286641417567
C_1_76 n447 PAR_2_1_VSS 9.82166251613e-11
R_2_76 PAR_0_2_VSS n448 0.633889059424
C_2_76 n448 PAR_2_1_VSS 2.84766445808e-10
R_3_76 PAR_0_2_VSS n449 0.85167468678
C_3_76 n449 PAR_2_1_VSS 4.42602189103e-10
R_4_76 PAR_0_2_VSS n450 1.94972128832
C_4_76 n450 PAR_2_1_VSS 4.9458858678e-10
R_5_76 PAR_0_2_VSS n451 3.55662698003
C_5_76 n451 PAR_2_1_VSS 1.14446575635e-09
R_6_76 PAR_0_2_VSS n452 9.72575139314
C_6_76 n452 PAR_2_1_VSS 1.41340132324e-09
G0_77 PAR_0_2_VSS PAR_2_1_VDD075CPU PAR_0_2_VSS PAR_2_1_VDD075CPU -0.228350242063
C0_77 PAR_0_2_VSS PAR_2_1_VDD075CPU 1.45822484258e-10
R_1_77 PAR_0_2_VSS n453 0.239160000825
C_1_77 n453 PAR_2_1_VDD075CPU 8.75760017339e-11
R_2_77 PAR_0_2_VSS n454 0.431556932141
C_2_77 n454 PAR_2_1_VDD075CPU 1.98638588837e-10
L_3_77 PAR_0_2_VSS n455 1.59373328125e-09
R_3_77 n455 PAR_2_1_VDD075CPU 4.72638281239
L_4_77 PAR_0_2_VSS n456 9.55934460969e-08
R_4_77 n456 PAR_2_1_VDD075CPU 59.6233469971
R_5_77 PAR_0_2_VSS n457 24.5374454314
C_5_77 n457 PAR_2_1_VDD075CPU 2.98451645697e-10
R0_78 PAR_0_2_VSS PAR_0_0_VSS 0.23107087874
C0_78 PAR_0_2_VSS PAR_0_0_VSS 2.15802306548e-10
R_1_78 PAR_0_2_VSS n458 0.0297793495978
C_1_78 n458 PAR_0_0_VSS 1.23225206064e-09
R_2_78 PAR_0_2_VSS n459 0.0551621452152
C_2_78 n459 PAR_0_0_VSS 2.27459570837e-09
R_3_78 PAR_0_2_VSS n460 0.078894209704
C_3_78 n460 PAR_0_0_VSS 3.63868623353e-09
R_4_78 PAR_0_2_VSS n461 0.158006543371
C_4_78 n461 PAR_0_0_VSS 6.5335027436e-09
R_5_78 PAR_0_2_VSS n462 0.402804982679
C_5_78 n462 PAR_0_0_VSS 9.202196097e-09
R_6_78 PAR_0_2_VSS n463 0.973230488495
C_6_78 n463 PAR_0_0_VSS 1.47568870231e-08
G0_79 PAR_0_2_VDD075CPU PAR_0_0_VDD075CPU PAR_0_2_VDD075CPU PAR_0_0_VDD075CPU -6.77933726032
C0_79 PAR_0_2_VDD075CPU PAR_0_0_VDD075CPU 1.30362353916e-10
R_1_79 PAR_0_2_VDD075CPU n464 0.394991094025
C_1_79 n464 PAR_0_0_VDD075CPU 7.47290325691e-11
L_2_79 PAR_0_2_VDD075CPU n465 1.7419146971e-11
R_2_79 n465 PAR_0_0_VDD075CPU 0.177891547402
R_3_79 PAR_0_2_VDD075CPU n466 0.265418229724
C_3_79 n466 PAR_0_0_VDD075CPU 5.33632301508e-10
L_4_79 PAR_0_2_VDD075CPU n467 3.88492310809e-10
R_4_79 n467 PAR_0_0_VDD075CPU 1.00388207433
R_5_79 PAR_0_2_VDD075CPU n468 2.19827000607
C_5_79 n468 PAR_0_0_VDD075CPU 4.22689439566e-10
L_6_79 PAR_0_2_VDD075CPU n469 1.93591243462e-08
R_6_79 n469 PAR_0_0_VDD075CPU 6.18222751636
R_7_79 PAR_0_2_VDD075CPU n470 39.8522061056
C_7_79 n470 PAR_0_0_VDD075CPU 3.31927856568e-10
G0_80 PAR_0_2_VDD075CPU PAR_1_0_VSS PAR_0_2_VDD075CPU PAR_1_0_VSS -0.491026640593
C0_80 PAR_0_2_VDD075CPU PAR_1_0_VSS 1.88987413731e-10
R_1_80 PAR_0_2_VDD075CPU n471 0.236576146158
C_1_80 n471 PAR_1_0_VSS 1.058286348e-10
R_2_80 PAR_0_2_VDD075CPU n472 0.705147361415
C_2_80 n472 PAR_1_0_VSS 1.45011649336e-10
L_3_80 PAR_0_2_VDD075CPU n473 7.20776221577e-10
R_3_80 n473 PAR_1_0_VSS 2.4810631744
L_4_80 PAR_0_2_VDD075CPU n474 2.17373022978e-08
R_4_80 n474 PAR_1_0_VSS 13.1946595458
L_5_80 PAR_0_2_VDD075CPU n475 8.20818679856e-07
R_5_80 n475 PAR_1_0_VSS 82.0655095927
G0_81 PAR_0_2_VDD075CPU PAR_1_0_VDD075CPU PAR_0_2_VDD075CPU PAR_1_0_VDD075CPU -3.73338293258
C0_81 PAR_0_2_VDD075CPU PAR_1_0_VDD075CPU 1.43433785254e-10
R_1_81 PAR_0_2_VDD075CPU n476 0.339522503539
C_1_81 n476 PAR_1_0_VDD075CPU 6.1160964518e-11
L_2_81 PAR_0_2_VDD075CPU n477 1.80411614026e-11
R_2_81 n477 PAR_1_0_VDD075CPU 0.313925901317
R_3_81 PAR_0_2_VDD075CPU n478 1.70171707213
C_3_81 n478 PAR_1_0_VDD075CPU 7.03514850075e-11
L_4_81 PAR_0_2_VDD075CPU n479 6.08648563081e-10
R_4_81 n479 PAR_1_0_VDD075CPU 2.08125565243
R_5_81 PAR_0_2_VDD075CPU n480 5.26373150389
C_5_81 n480 PAR_1_0_VDD075CPU 1.2743608227e-10
L_6_81 PAR_0_2_VDD075CPU n481 3.5257584972e-08
R_6_81 n481 PAR_1_0_VDD075CPU 15.3366954397
R_7_81 PAR_0_2_VDD075CPU n482 95.7028042311
C_7_81 n482 PAR_1_0_VDD075CPU 1.20769490879e-10
L_8_81 PAR_0_2_VDD075CPU n483 0.0155329587949
R_8_81 n483 PAR_1_0_VDD075CPU 425.772987646
G0_82 PAR_0_2_VDD075CPU PAR_2_0_VSS PAR_0_2_VDD075CPU PAR_2_0_VSS -0.117529860111
C0_82 PAR_0_2_VDD075CPU PAR_2_0_VSS 2.19380010451e-10
R_1_82 PAR_0_2_VDD075CPU n484 3.37550910325
C_1_82 n484 PAR_2_0_VSS 1.24991072667e-11
R_2_82 PAR_0_2_VDD075CPU n485 4.52065134713
C_2_82 n485 PAR_2_0_VSS 2.9104364337e-11
R_3_82 PAR_0_2_VDD075CPU n486 4.72197110057
C_3_82 n486 PAR_2_0_VSS 1.20793943171e-10
L_4_82 PAR_0_2_VDD075CPU n487 1.58544204195e-08
R_4_82 n487 PAR_2_0_VSS 10.3478274529
L_5_82 PAR_0_2_VDD075CPU n488 3.31211232174e-07
R_5_82 n488 PAR_2_0_VSS 69.7768997738
L_6_82 PAR_0_2_VDD075CPU n489 2.26982633849e-06
R_6_82 n489 PAR_2_0_VSS 152.442986826
G0_83 PAR_0_2_VDD075CPU PAR_2_0_VDD075CPU PAR_0_2_VDD075CPU PAR_2_0_VDD075CPU -3.79676078189
C0_83 PAR_0_2_VDD075CPU PAR_2_0_VDD075CPU 1.56009061894e-10
R_1_83 PAR_0_2_VDD075CPU n490 0.319441915483
C_1_83 n490 PAR_2_0_VDD075CPU 6.61117680118e-11
L_2_83 PAR_0_2_VDD075CPU n491 1.70935985154e-11
R_2_83 n491 PAR_2_0_VDD075CPU 0.306242625973
R_3_83 PAR_0_2_VDD075CPU n492 2.08339822011
C_3_83 n492 PAR_2_0_VDD075CPU 5.9292851591e-11
L_4_83 PAR_0_2_VDD075CPU n493 6.49430149493e-10
R_4_83 n493 PAR_2_0_VDD075CPU 2.12626385193
R_5_83 PAR_0_2_VDD075CPU n494 5.59548440299
C_5_83 n494 PAR_2_0_VDD075CPU 1.24638134251e-10
L_6_83 PAR_0_2_VDD075CPU n495 4.13281488732e-08
R_6_83 n495 PAR_2_0_VDD075CPU 16.3983921909
R_7_83 PAR_0_2_VDD075CPU n496 131.568064579
C_7_83 n496 PAR_2_0_VDD075CPU 9.2362203906e-11
G0_84 PAR_0_2_VDD075CPU PAR_0_1_VSS PAR_0_2_VDD075CPU PAR_0_1_VSS -0.0342870164517
C0_84 PAR_0_2_VDD075CPU PAR_0_1_VSS 1.79198548429e-10
R_1_84 PAR_0_2_VDD075CPU n497 0.0527145214051
C_1_84 n497 PAR_0_1_VSS 2.71068993508e-10
R_2_84 PAR_0_2_VDD075CPU n498 0.106475709056
C_2_84 n498 PAR_0_1_VSS 4.36401058396e-10
R_3_84 PAR_0_2_VDD075CPU n499 0.0228553105165
C_3_84 n499 PAR_0_1_VSS 4.43301205782e-09
L_4_84 PAR_0_2_VDD075CPU n500 1.53863404329e-08
R_4_84 n500 PAR_0_1_VSS 29.1655566291
R_5_84 PAR_0_2_VDD075CPU n501 26.9281278009
C_5_84 n501 PAR_0_1_VSS 1.52684524497e-10
R_6_84 PAR_0_2_VDD075CPU n502 54.8376001505
C_6_84 n502 PAR_0_1_VSS 2.56319452408e-10
R0_85 PAR_0_2_VDD075CPU PAR_0_1_VDD075CPU 0.00586625090786
C0_85 PAR_0_2_VDD075CPU PAR_0_1_VDD075CPU 4.75556803258e-11
L_1_85 PAR_0_2_VDD075CPU n503 1.43305506522e-12
R_1_85 n503 PAR_0_1_VDD075CPU 0.0925128490814
L_2_85 PAR_0_2_VDD075CPU n504 9.25890016161e-12
R_2_85 n504 PAR_0_1_VDD075CPU 0.195013544553
L_3_85 PAR_0_2_VDD075CPU n505 3.47360740477e-12
R_3_85 n505 PAR_0_1_VDD075CPU 0.0337850258666
L_4_85 PAR_0_2_VDD075CPU n506 2.23782833039e-08
R_4_85 n506 PAR_0_1_VDD075CPU 45.6913978982
L_5_85 PAR_0_2_VDD075CPU n507 1.40124615801e-06
R_5_85 n507 PAR_0_1_VDD075CPU 441.586210734
G0_86 PAR_0_2_VDD075CPU PAR_1_1_VSS PAR_0_2_VDD075CPU PAR_1_1_VSS -2.23878071967
C0_86 PAR_0_2_VDD075CPU PAR_1_1_VSS 9.96187252199e-11
R_1_86 PAR_0_2_VDD075CPU n508 2.27531929011
C_1_86 n508 PAR_1_1_VSS 6.90619304127e-12
L_2_86 PAR_0_2_VDD075CPU n509 2.50231730847e-11
R_2_86 n509 PAR_1_1_VSS 0.538410127986
R_3_86 PAR_0_2_VDD075CPU n510 0.589542018573
C_3_86 n510 PAR_1_1_VSS 1.76619322125e-10
L_4_86 PAR_0_2_VDD075CPU n511 5.60895671017e-10
R_4_86 n511 PAR_1_1_VSS 2.98710763971
R_5_86 PAR_0_2_VDD075CPU n512 10.8984398867
C_5_86 n512 PAR_1_1_VSS 4.04788774953e-11
L_6_86 PAR_0_2_VDD075CPU n513 2.5048336626e-08
R_6_86 n513 PAR_1_1_VSS 23.1995394404
R_7_86 PAR_0_2_VDD075CPU n514 88.5443651526
C_7_86 n514 PAR_1_1_VSS 3.94355634876e-11
L_8_86 PAR_0_2_VDD075CPU n515 3.84087877832e-06
R_8_86 n515 PAR_1_1_VSS 278.999957249
R0_87 PAR_0_2_VDD075CPU PAR_1_1_VDD075CPU 0.33715892405
C0_87 PAR_0_2_VDD075CPU PAR_1_1_VDD075CPU 1.23417458362e-10
L_1_87 PAR_0_2_VDD075CPU n516 5.06001696106e-12
R_1_87 n516 PAR_1_1_VDD075CPU 0.286783632071
L_2_87 PAR_0_2_VDD075CPU n517 9.25784964039e-11
R_2_87 n517 PAR_1_1_VDD075CPU 1.53985643633
L_3_87 PAR_0_2_VDD075CPU n518 6.13317153798e-11
R_3_87 n518 PAR_1_1_VDD075CPU 0.569361217875
L_4_87 PAR_0_2_VDD075CPU n519 2.10035492123e-08
R_4_87 n519 PAR_1_1_VDD075CPU 52.6634597533
L_5_87 PAR_0_2_VDD075CPU n520 5.07653336955e-07
R_5_87 n520 PAR_1_1_VDD075CPU 345.616257927
L_6_87 PAR_0_2_VDD075CPU n521 2.17661602436e-05
R_6_87 n521 PAR_1_1_VDD075CPU 1919.75424607
G0_88 PAR_0_2_VDD075CPU PAR_2_1_VSS PAR_0_2_VDD075CPU PAR_2_1_VSS -1.32324939607
C0_88 PAR_0_2_VDD075CPU PAR_2_1_VSS 1.25282210633e-10
R_1_88 PAR_0_2_VDD075CPU n522 1.60662970664
C_1_88 n522 PAR_2_1_VSS 1.36746557552e-11
L_2_88 PAR_0_2_VDD075CPU n523 1.0044650193e-10
R_2_88 n523 PAR_2_1_VSS 1.20030165659
R_3_88 PAR_0_2_VDD075CPU n524 2.09024201716
C_3_88 n524 PAR_2_1_VSS 1.07706273744e-10
L_4_88 PAR_0_2_VDD075CPU n525 1.45944835165e-09
R_4_88 n525 PAR_2_1_VSS 2.57046295595
R_5_88 PAR_0_2_VDD075CPU n526 4.83271890741
C_5_88 n526 PAR_2_1_VSS 2.98040921352e-10
L_6_88 PAR_0_2_VDD075CPU n527 4.13185179606e-08
R_6_88 n527 PAR_2_1_VSS 9.89212457502
R_7_88 PAR_0_2_VDD075CPU n528 64.549102582
C_7_88 n528 PAR_2_1_VSS 2.20636232668e-10
G0_89 PAR_0_2_VDD075CPU PAR_2_1_VDD075CPU PAR_0_2_VDD075CPU PAR_2_1_VDD075CPU -2.45970019813
C0_89 PAR_0_2_VDD075CPU PAR_2_1_VDD075CPU 1.07566999834e-10
R_1_89 PAR_0_2_VDD075CPU n529 0.434205783279
C_1_89 n529 PAR_2_1_VDD075CPU 4.98803282939e-11
L_2_89 PAR_0_2_VDD075CPU n530 2.34191000329e-11
R_2_89 n530 PAR_2_1_VDD075CPU 0.453244136065
R_3_89 PAR_0_2_VDD075CPU n531 20.1116571989
C_3_89 n531 PAR_2_1_VDD075CPU 6.19374135268e-12
L_4_89 PAR_0_2_VDD075CPU n532 1.78314584372e-09
R_4_89 n532 PAR_2_1_VDD075CPU 4.81344984693
R_5_89 PAR_0_2_VDD075CPU n533 10.1892099555
C_5_89 n533 PAR_2_1_VDD075CPU 9.22746103862e-11
L_6_89 PAR_0_2_VDD075CPU n534 7.20903317184e-08
R_6_89 n534 PAR_2_1_VDD075CPU 22.7596971237
R_7_89 PAR_0_2_VDD075CPU n535 113.904360169
C_7_89 n535 PAR_2_1_VDD075CPU 1.17057027714e-10
L_8_89 PAR_0_2_VDD075CPU n536 0.0243497818825
R_8_89 n536 PAR_2_1_VDD075CPU 542.866832645
C0_90 PAR_0_2_VDD075CPU PAR_0_2_VSS 2.25484535946e-10
R_1_90 PAR_0_2_VDD075CPU n537 0.00144166038323
C_1_90 n537 PAR_0_2_VSS 1.39076681527e-08
R_2_90 PAR_0_2_VDD075CPU n538 0.000819926062675
C_2_90 n538 PAR_0_2_VSS 4.73783009406e-08
R_3_90 PAR_0_2_VDD075CPU n539 0.00356045721808
C_3_90 n539 PAR_0_2_VSS 2.71451909962e-08
R_4_90 PAR_0_2_VDD075CPU n540 0.820914742475
C_4_90 n540 PAR_0_2_VSS 3.35661239235e-10
R_5_90 PAR_0_2_VDD075CPU n541 12.4149966998
C_5_90 n541 PAR_0_2_VSS 9.45028414109e-11
R_6_90 PAR_0_2_VDD075CPU n542 23.7226630167
C_6_90 n542 PAR_0_2_VSS 3.44822442363e-10
G0_91 PAR_0_2_VDD075CPU PAR_0_0_VSS PAR_0_2_VDD075CPU PAR_0_0_VSS -0.934406822118
C0_91 PAR_0_2_VDD075CPU PAR_0_0_VSS 2.31279955209e-10
R_1_91 PAR_0_2_VDD075CPU n543 0.0171143553403
C_1_91 n543 PAR_0_0_VSS 8.61217060097e-10
R_2_91 PAR_0_2_VDD075CPU n544 0.8697663411
C_2_91 n544 PAR_0_0_VSS 7.12827650003e-11
L_3_91 PAR_0_2_VDD075CPU n545 2.52530822661e-10
R_3_91 n545 PAR_0_0_VSS 1.07019766269
R_4_91 PAR_0_2_VDD075CPU n546 14.173192481
C_4_91 n546 PAR_0_0_VSS 8.09649622756e-11
R_5_91 PAR_0_2_VDD075CPU n547 87.7703323089
C_5_91 n547 PAR_0_0_VSS 1.07029649908e-10
G0_92 PAR_1_2_VSS PAR_0_0_VDD075CPU PAR_1_2_VSS PAR_0_0_VDD075CPU -0.803101940207
C0_92 PAR_1_2_VSS PAR_0_0_VDD075CPU 1.43445191696e-10
R_1_92 PAR_1_2_VSS n548 0.115511116085
C_1_92 n548 PAR_0_0_VDD075CPU 4.85382260503e-11
R_2_92 PAR_1_2_VSS n549 1.01243352442
C_2_92 n549 PAR_0_0_VDD075CPU 5.23240167911e-11
R_3_92 PAR_1_2_VSS n550 1.51407937859
C_3_92 n550 PAR_0_0_VDD075CPU 1.09242515486e-10
L_4_92 PAR_1_2_VSS n551 2.34551645698e-10
R_4_92 n551 PAR_0_0_VDD075CPU 1.28670160925
R_5_92 PAR_1_2_VSS n552 17.4276302497
C_5_92 n552 PAR_0_0_VDD075CPU 3.79449564719e-11
L_6_92 PAR_1_2_VSS n553 2.26607147649e-07
R_6_92 n553 PAR_0_0_VDD075CPU 54.381381661
L_7_92 PAR_1_2_VSS n554 1.87684789413e-06
R_7_92 n554 PAR_0_0_VDD075CPU 132.761050956
G0_93 PAR_1_2_VSS PAR_1_0_VSS PAR_1_2_VSS PAR_1_0_VSS -0.339375632033
C0_93 PAR_1_2_VSS PAR_1_0_VSS 1.70007521837e-10
R_1_93 PAR_1_2_VSS n555 0.327756461696
C_1_93 n555 PAR_1_0_VSS 1.347315529e-10
R_2_93 PAR_1_2_VSS n556 0.703273412338
C_2_93 n556 PAR_1_0_VSS 2.01951623041e-10
R_3_93 PAR_1_2_VSS n557 0.347569853095
C_3_93 n557 PAR_1_0_VSS 6.45896512378e-10
R_4_93 PAR_1_2_VSS n558 0.37772974527
C_4_93 n558 PAR_1_0_VSS 2.64064701706e-09
L_5_93 PAR_1_2_VSS n559 2.11552197763e-08
R_5_93 n559 PAR_1_0_VSS 4.09164695662
L_6_93 PAR_1_2_VSS n560 1.6088458232e-07
R_6_93 n560 PAR_1_0_VSS 10.5290467836
G0_94 PAR_1_2_VSS PAR_1_0_VDD075CPU PAR_1_2_VSS PAR_1_0_VDD075CPU -0.228233462774
C0_94 PAR_1_2_VSS PAR_1_0_VDD075CPU 1.77394909501e-10
R_1_94 PAR_1_2_VSS n561 0.842800648578
C_1_94 n561 PAR_1_0_VDD075CPU 5.48121910444e-11
R_2_94 PAR_1_2_VSS n562 3.28551555423
C_2_94 n562 PAR_1_0_VDD075CPU 3.05816908748e-11
L_3_94 PAR_1_2_VSS n563 1.03612573009e-09
R_3_94 n563 PAR_1_0_VDD075CPU 4.89268704261
R_4_94 PAR_1_2_VSS n564 16.3334510499
C_4_94 n564 PAR_1_0_VDD075CPU 4.18329618461e-11
L_5_94 PAR_1_2_VSS n565 2.92528171848e-07
R_5_94 n565 PAR_1_0_VDD075CPU 59.1806700585
L_6_94 PAR_1_2_VSS n566 2.16493405066e-06
R_6_94 n566 PAR_1_0_VDD075CPU 143.897558561
G0_95 PAR_1_2_VSS PAR_2_0_VSS PAR_1_2_VSS PAR_2_0_VSS -0.798517718533
C0_95 PAR_1_2_VSS PAR_2_0_VSS 1.98754002106e-10
R_1_95 PAR_1_2_VSS n567 0.46333512947
C_1_95 n567 PAR_2_0_VSS 1.00901285275e-10
R_2_95 PAR_1_2_VSS n568 1.05259000686
C_2_95 n568 PAR_2_0_VSS 1.62478385363e-10
R_3_95 PAR_1_2_VSS n569 0.257466274123
C_3_95 n569 PAR_2_0_VSS 4.50114487319e-09
L_4_95 PAR_1_2_VSS n570 4.28327992794e-09
R_4_95 n570 PAR_2_0_VSS 1.65771181904
L_5_95 PAR_1_2_VSS n571 5.93903121779e-08
R_5_95 n571 PAR_2_0_VSS 5.12094149951
G0_96 PAR_1_2_VSS PAR_2_0_VDD075CPU PAR_1_2_VSS PAR_2_0_VDD075CPU -0.036786241754
C0_96 PAR_1_2_VSS PAR_2_0_VDD075CPU 1.92345065599e-10
R_1_96 PAR_1_2_VSS n572 0.694482157719
C_1_96 n572 PAR_2_0_VDD075CPU 7.9143060805e-11
R_2_96 PAR_1_2_VSS n573 19.3657808419
C_2_96 n573 PAR_2_0_VDD075CPU 5.9486369148e-11
L_3_96 PAR_1_2_VSS n574 1.44736455499e-07
R_3_96 n574 PAR_2_0_VDD075CPU 27.1840745869
R0_97 PAR_1_2_VSS PAR_0_1_VSS 0.123785961561
C0_97 PAR_1_2_VSS PAR_0_1_VSS 1.60127311906e-10
R_1_97 PAR_1_2_VSS n575 0.278064437794
C_1_97 n575 PAR_0_1_VSS 1.75787138906e-10
R_2_97 PAR_1_2_VSS n576 0.326834215634
C_2_97 n576 PAR_0_1_VSS 5.37801629899e-10
R_3_97 PAR_1_2_VSS n577 0.659470146978
C_3_97 n577 PAR_0_1_VSS 5.70511615393e-10
R_4_97 PAR_1_2_VSS n578 0.558307551107
C_4_97 n578 PAR_0_1_VSS 1.87933550215e-09
R_5_97 PAR_1_2_VSS n579 0.915535426194
C_5_97 n579 PAR_0_1_VSS 4.04525024307e-09
R_6_97 PAR_1_2_VSS n580 2.94963409779
C_6_97 n580 PAR_0_1_VSS 4.65501593935e-09
G0_98 PAR_1_2_VSS PAR_0_1_VDD075CPU PAR_1_2_VSS PAR_0_1_VDD075CPU -0.0275569743297
C0_98 PAR_1_2_VSS PAR_0_1_VDD075CPU 1.39028720157e-10
R_1_98 PAR_1_2_VSS n581 0.932344663353
C_1_98 n581 PAR_0_1_VDD075CPU 3.31284596363e-11
R_2_98 PAR_1_2_VSS n582 1.15491429906
C_2_98 n582 PAR_0_1_VDD075CPU 8.01785187582e-11
R_3_98 PAR_1_2_VSS n583 25.177362109
C_3_98 n583 PAR_0_1_VDD075CPU 5.27654641844e-11
L_4_98 PAR_1_2_VSS n584 1.96921294964e-07
R_4_98 n584 PAR_0_1_VDD075CPU 36.2884512653
R0_99 PAR_1_2_VSS PAR_1_1_VSS 0.00605155316325
C0_99 PAR_1_2_VSS PAR_1_1_VSS 7.52440640938e-12
L_1_99 PAR_1_2_VSS n585 1.95832559308e-12
R_1_99 n585 PAR_1_1_VSS 0.133342404264
L_2_99 PAR_1_2_VSS n586 1.55434810905e-10
R_2_99 n586 PAR_1_1_VSS 2.65479066948
L_3_99 PAR_1_2_VSS n587 5.59706832147e-12
R_3_99 n587 PAR_1_1_VSS 0.0538633214303
R_4_99 PAR_1_2_VSS n588 33.8661992693
C_4_99 n588 PAR_1_1_VSS 2.21834169607e-11
L_5_99 PAR_1_2_VSS n589 5.94821862127e-07
R_5_99 n589 PAR_1_1_VSS 118.397647693
L_6_99 PAR_1_2_VSS n590 4.78697622246e-06
R_6_99 n590 PAR_1_1_VSS 309.437645508
G0_100 PAR_1_2_VSS PAR_1_1_VDD075CPU PAR_1_2_VSS PAR_1_1_VDD075CPU -0.0150457184579
C0_100 PAR_1_2_VSS PAR_1_1_VDD075CPU 1.23183886518e-10
R_1_100 PAR_1_2_VSS n591 0.314945268321
C_1_100 n591 PAR_1_1_VDD075CPU 8.25887895379e-11
R_2_100 PAR_1_2_VSS n592 0.0753596989232
C_2_100 n592 PAR_1_1_VDD075CPU 1.39055193494e-09
R_3_100 PAR_1_2_VSS n593 28.2009607936
C_3_100 n593 PAR_1_1_VDD075CPU 3.28745574383e-11
L_4_100 PAR_1_2_VSS n594 4.52425230553e-07
R_4_100 n594 PAR_1_1_VDD075CPU 66.4640815086
R0_101 PAR_1_2_VSS PAR_2_1_VSS 1.7983778067
C0_101 PAR_1_2_VSS PAR_2_1_VSS 1.37366070454e-10
R_1_101 PAR_1_2_VSS n595 1.08239914123
C_1_101 n595 PAR_2_1_VSS 4.24378073427e-11
L_2_101 PAR_1_2_VSS n596 2.3610679026e-11
R_2_101 n596 PAR_2_1_VSS 0.156944433032
R_3_101 PAR_1_2_VSS n597 0.138579228034
C_3_101 n597 PAR_2_1_VSS 1.40070044462e-09
L_4_101 PAR_1_2_VSS n598 2.76338429306e-10
R_4_101 n598 PAR_2_1_VSS 0.448071301838
L_5_101 PAR_1_2_VSS n599 8.0790092772e-10
R_5_101 n599 PAR_2_1_VSS 0.6829495994
L_6_101 PAR_1_2_VSS n600 2.71782654199e-08
R_6_101 n600 PAR_2_1_VSS 6.86027617156
L_7_101 PAR_1_2_VSS n601 3.38140733381e-07
R_7_101 n601 PAR_2_1_VSS 24.0799472798
G0_102 PAR_1_2_VSS PAR_2_1_VDD075CPU PAR_1_2_VSS PAR_2_1_VDD075CPU -1.14462662796
C0_102 PAR_1_2_VSS PAR_2_1_VDD075CPU 1.30464562192e-10
R_1_102 PAR_1_2_VSS n602 1.18141304558
C_1_102 n602 PAR_2_1_VDD075CPU 3.58125715087e-11
R_2_102 PAR_1_2_VSS n603 0.493862406032
C_2_102 n603 PAR_2_1_VDD075CPU 2.72952461806e-10
L_3_102 PAR_1_2_VSS n604 1.66692213719e-10
R_3_102 n604 PAR_2_1_VDD075CPU 0.884086535856
R_4_102 PAR_1_2_VSS n605 7.241289978
C_4_102 n605 PAR_2_1_VDD075CPU 1.07198910744e-10
L_5_102 PAR_1_2_VSS n606 6.65273751669e-07
R_5_102 n606 PAR_2_1_VDD075CPU 73.9883760781
R0_103 PAR_1_2_VSS PAR_0_2_VSS 0.00387436069848
L_1_103 PAR_1_2_VSS n607 7.67628811718e-13
R_1_103 n607 PAR_0_2_VSS 0.0244601689327
L_2_103 PAR_1_2_VSS n608 7.39652813295e-12
R_2_103 n608 PAR_0_2_VSS 0.0799763682914
R_3_103 PAR_1_2_VSS n609 0.46967540487
C_3_103 n609 PAR_0_2_VSS 5.97261383511e-10
R_4_103 PAR_1_2_VSS n610 0.521500517726
C_4_103 n610 PAR_0_2_VSS 1.90506975718e-09
R_5_103 PAR_1_2_VSS n611 0.963456664776
C_5_103 n611 PAR_0_2_VSS 3.89330958558e-09
R_6_103 PAR_1_2_VSS n612 2.97575143829
C_6_103 n612 PAR_0_2_VSS 4.43567586768e-09
G0_104 PAR_1_2_VSS PAR_0_2_VDD075CPU PAR_1_2_VSS PAR_0_2_VDD075CPU -0.021596066111
C0_104 PAR_1_2_VSS PAR_0_2_VDD075CPU 1.68979660067e-10
R_1_104 PAR_1_2_VSS n613 0.0342399022335
C_1_104 n613 PAR_0_2_VDD075CPU 1.01070758482e-09
R_2_104 PAR_1_2_VSS n614 0.0917877582928
C_2_104 n614 PAR_0_2_VDD075CPU 1.09621677288e-09
R_3_104 PAR_1_2_VSS n615 42.718002961
C_3_104 n615 PAR_0_2_VDD075CPU 3.45351658031e-11
L_4_104 PAR_1_2_VSS n616 4.02931030026e-07
R_4_104 n616 PAR_0_2_VDD075CPU 46.3047246095
R0_105 PAR_1_2_VSS PAR_0_0_VSS 47929.1493764
C0_105 PAR_1_2_VSS PAR_0_0_VSS 2.6561331623e-10
R_1_105 PAR_1_2_VSS n617 0.0365201730577
C_1_105 n617 PAR_0_0_VSS 7.31845820601e-10
R_2_105 PAR_1_2_VSS n618 0.119756969806
C_2_105 n618 PAR_0_0_VSS 6.77311876519e-10
R_3_105 PAR_1_2_VSS n619 0.165514575802
C_3_105 n619 PAR_0_0_VSS 1.28360029738e-09
R_4_105 PAR_1_2_VSS n620 0.208579023405
C_4_105 n620 PAR_0_0_VSS 5.49679069501e-09
R_5_105 PAR_1_2_VSS n621 0.331075847408
C_5_105 n621 PAR_0_0_VSS 7.38616550371e-09
R_6_105 PAR_1_2_VSS n622 6.21643858683
C_6_105 n622 PAR_0_0_VSS 1.87101928604e-09
G0_106 PAR_1_2_VDD075CPU PAR_0_0_VDD075CPU PAR_1_2_VDD075CPU PAR_0_0_VDD075CPU -4.95010367129
C0_106 PAR_1_2_VDD075CPU PAR_0_0_VDD075CPU 1.27022794937e-10
R_1_106 PAR_1_2_VDD075CPU n623 0.37048143233
C_1_106 n623 PAR_0_0_VDD075CPU 6.85789698024e-11
L_2_106 PAR_1_2_VDD075CPU n624 1.84794633188e-11
R_2_106 n624 PAR_0_0_VDD075CPU 0.242209821857
R_3_106 PAR_1_2_VDD075CPU n625 0.524185834121
C_3_106 n625 PAR_0_0_VDD075CPU 2.49848592521e-10
L_4_106 PAR_1_2_VDD075CPU n626 5.14441066062e-10
R_4_106 n626 PAR_0_0_VDD075CPU 1.42253076263
R_5_106 PAR_1_2_VDD075CPU n627 3.06073806438
C_5_106 n627 PAR_0_0_VDD075CPU 2.82278101524e-10
L_6_106 PAR_1_2_VDD075CPU n628 2.43881249845e-08
R_6_106 n628 PAR_0_0_VDD075CPU 8.42659611737
R_7_106 PAR_1_2_VDD075CPU n629 60.7013219838
C_7_106 n629 PAR_0_0_VDD075CPU 2.14310704887e-10
G0_107 PAR_1_2_VDD075CPU PAR_1_0_VSS PAR_1_2_VDD075CPU PAR_1_0_VSS -0.313926047527
C0_107 PAR_1_2_VDD075CPU PAR_1_0_VSS 1.93620677266e-10
R_1_107 PAR_1_2_VDD075CPU n630 0.322643245386
C_1_107 n630 PAR_1_0_VSS 8.2198410627e-11
R_2_107 PAR_1_2_VDD075CPU n631 0.974668548479
C_2_107 n631 PAR_1_0_VSS 1.16323106203e-10
L_3_107 PAR_1_2_VDD075CPU n632 1.32330693991e-09
R_3_107 n632 PAR_1_0_VSS 4.35153029924
L_4_107 PAR_1_2_VDD075CPU n633 2.37506158896e-08
R_4_107 n633 PAR_1_0_VSS 13.7016741557
L_5_107 PAR_1_2_VDD075CPU n634 9.60363137532e-07
R_5_107 n634 PAR_1_0_VSS 89.7822940015
G0_108 PAR_1_2_VDD075CPU PAR_1_0_VDD075CPU PAR_1_2_VDD075CPU PAR_1_0_VDD075CPU -4.24419613475
C0_108 PAR_1_2_VDD075CPU PAR_1_0_VDD075CPU 1.40244845484e-10
R_1_108 PAR_1_2_VDD075CPU n635 0.334523451799
C_1_108 n635 PAR_1_0_VDD075CPU 5.0013179453e-11
L_2_108 PAR_1_2_VDD075CPU n636 1.56589997741e-11
R_2_108 n636 PAR_1_0_VDD075CPU 0.300927501523
R_3_108 PAR_1_2_VDD075CPU n637 1.10667379438
C_3_108 n637 PAR_1_0_VDD075CPU 1.06385649573e-10
L_4_108 PAR_1_2_VDD075CPU n638 3.04108813608e-10
R_4_108 n638 PAR_1_0_VDD075CPU 1.31624206721
R_5_108 PAR_1_2_VDD075CPU n639 3.24494705077
C_5_108 n639 PAR_1_0_VDD075CPU 1.62350263306e-10
L_6_108 PAR_1_2_VDD075CPU n640 8.37044197516e-09
R_6_108 n640 PAR_1_0_VDD075CPU 6.70517227313
R_7_108 PAR_1_2_VDD075CPU n641 23.2077693463
C_7_108 n641 PAR_1_0_VDD075CPU 1.63946176004e-10
L_8_108 PAR_1_2_VDD075CPU n642 1.16107801352e-06
R_8_108 n642 PAR_1_0_VDD075CPU 82.3826987677
G0_109 PAR_1_2_VDD075CPU PAR_2_0_VSS PAR_1_2_VDD075CPU PAR_2_0_VSS -0.427096170162
C0_109 PAR_1_2_VDD075CPU PAR_2_0_VSS 2.11314823748e-10
L_1_109 PAR_1_2_VDD075CPU n643 2.08221295285e-11
R_1_109 n643 PAR_2_0_VSS 3.23610614916
R_2_109 PAR_1_2_VDD075CPU n644 6.7453502733
C_2_109 n644 PAR_2_0_VSS 2.25394375135e-11
R_3_109 PAR_1_2_VDD075CPU n645 3.58621016057
C_3_109 n645 PAR_2_0_VSS 1.50394598284e-10
L_4_109 PAR_1_2_VDD075CPU n646 1.68278889814e-08
R_4_109 n646 PAR_2_0_VSS 9.22465999044
L_5_109 PAR_1_2_VDD075CPU n647 1.13770122335e-06
R_5_109 n647 PAR_2_0_VSS 103.329873557
G0_110 PAR_1_2_VDD075CPU PAR_2_0_VDD075CPU PAR_1_2_VDD075CPU PAR_2_0_VDD075CPU -4.33552628806
C0_110 PAR_1_2_VDD075CPU PAR_2_0_VDD075CPU 1.52203946349e-10
R_1_110 PAR_1_2_VDD075CPU n648 0.321818809581
C_1_110 n648 PAR_2_0_VDD075CPU 5.22086633137e-11
L_2_110 PAR_1_2_VDD075CPU n649 1.52991410181e-11
R_2_110 n649 PAR_2_0_VDD075CPU 0.297805704929
R_3_110 PAR_1_2_VDD075CPU n650 1.26939960571
C_3_110 n650 PAR_2_0_VDD075CPU 9.62683553517e-11
L_4_110 PAR_1_2_VDD075CPU n651 3.26120583839e-10
R_4_110 n651 PAR_2_0_VDD075CPU 1.28325316355
R_5_110 PAR_1_2_VDD075CPU n652 2.54480661348
C_5_110 n652 PAR_2_0_VDD075CPU 2.09069083102e-10
L_6_110 PAR_1_2_VDD075CPU n653 6.36947857632e-09
R_6_110 n653 PAR_2_0_VDD075CPU 5.39656950776
R_7_110 PAR_1_2_VDD075CPU n654 21.0719056735
C_7_110 n654 PAR_2_0_VDD075CPU 1.71595639687e-10
L_8_110 PAR_1_2_VDD075CPU n655 1.05788761458e-06
R_8_110 n655 PAR_2_0_VDD075CPU 76.838857278
G0_111 PAR_1_2_VDD075CPU PAR_0_1_VSS PAR_1_2_VDD075CPU PAR_0_1_VSS -0.09734685759
C0_111 PAR_1_2_VDD075CPU PAR_0_1_VSS 1.9758971558e-10
R_1_111 PAR_1_2_VDD075CPU n656 0.155049263877
C_1_111 n656 PAR_0_1_VSS 1.66538199447e-10
R_2_111 PAR_1_2_VDD075CPU n657 0.217554864944
C_2_111 n657 PAR_0_1_VSS 4.58741377484e-10
L_3_111 PAR_1_2_VDD075CPU n658 5.91831308194e-09
R_3_111 n658 PAR_0_1_VSS 10.27254502
R_4_111 PAR_1_2_VDD075CPU n659 29.7075446916
C_4_111 n659 PAR_0_1_VSS 1.84526140988e-10
R_5_111 PAR_1_2_VDD075CPU n660 81.3464961603
C_5_111 n660 PAR_0_1_VSS 2.07635510528e-10
R0_112 PAR_1_2_VDD075CPU PAR_0_1_VDD075CPU 0.336621295623
C0_112 PAR_1_2_VDD075CPU PAR_0_1_VDD075CPU 1.48035883098e-10
L_1_112 PAR_1_2_VDD075CPU n661 5.97713499834e-12
R_1_112 n661 PAR_0_1_VDD075CPU 0.283732843103
L_2_112 PAR_1_2_VDD075CPU n662 7.17396524338e-11
R_2_112 n662 PAR_0_1_VDD075CPU 0.897715876079
L_3_112 PAR_1_2_VDD075CPU n663 8.38542869879e-11
R_3_112 n663 PAR_0_1_VDD075CPU 0.705699591856
L_4_112 PAR_1_2_VDD075CPU n664 2.40381799303e-08
R_4_112 n664 PAR_0_1_VDD075CPU 47.2592283588
L_5_112 PAR_1_2_VDD075CPU n665 1.19728425648e-06
R_5_112 n665 PAR_0_1_VDD075CPU 410.04468114
L_6_112 PAR_1_2_VDD075CPU n666 0.000469352105924
R_6_112 n666 PAR_0_1_VDD075CPU 2784.53707916
G0_113 PAR_1_2_VDD075CPU PAR_1_1_VSS PAR_1_2_VDD075CPU PAR_1_1_VSS -0.0176446748112
C0_113 PAR_1_2_VDD075CPU PAR_1_1_VSS 1.42450891029e-10
R_1_113 PAR_1_2_VDD075CPU n667 0.0764479016671
C_1_113 n667 PAR_1_1_VSS 1.51441314031e-10
R_2_113 PAR_1_2_VDD075CPU n668 0.128387654401
C_2_113 n668 PAR_1_1_VSS 3.94319976916e-10
R_3_113 PAR_1_2_VDD075CPU n669 0.0291237816826
C_3_113 n669 PAR_1_1_VSS 3.44101929275e-09
L_4_113 PAR_1_2_VDD075CPU n670 2.74557964147e-08
R_4_113 n670 PAR_1_1_VSS 67.7675514418
L_5_113 PAR_1_2_VDD075CPU n671 5.64320378101e-07
R_5_113 n671 PAR_1_1_VSS 407.611974853
L_6_113 PAR_1_2_VDD075CPU n672 2.2210747811e-05
R_6_113 n672 PAR_1_1_VSS 2298.6478252
R0_114 PAR_1_2_VDD075CPU PAR_1_1_VDD075CPU 0.0057171066167
C0_114 PAR_1_2_VDD075CPU PAR_1_1_VDD075CPU 3.05655419297e-11
L_1_114 PAR_1_2_VDD075CPU n673 8.42375582558e-13
R_1_114 n673 PAR_1_1_VDD075CPU 0.064323400611
L_2_114 PAR_1_2_VDD075CPU n674 8.29701718622e-12
R_2_114 n674 PAR_1_1_VDD075CPU 0.169995773317
L_3_114 PAR_1_2_VDD075CPU n675 3.95691376681e-12
R_3_114 n675 PAR_1_1_VDD075CPU 0.0388696104919
L_4_114 PAR_1_2_VDD075CPU n676 2.30291202994e-08
R_4_114 n676 PAR_1_1_VDD075CPU 53.3046290106
L_5_114 PAR_1_2_VDD075CPU n677 7.03110494024e-07
R_5_114 n677 PAR_1_1_VDD075CPU 381.719003272
L_6_114 PAR_1_2_VDD075CPU n678 9.62100124426e-05
R_6_114 n678 PAR_1_1_VDD075CPU 4875.33613937
G0_115 PAR_1_2_VDD075CPU PAR_2_1_VSS PAR_1_2_VDD075CPU PAR_2_1_VSS -5.51332987274
C0_115 PAR_1_2_VDD075CPU PAR_2_1_VSS 1.57325533589e-10
L_1_115 PAR_1_2_VDD075CPU n679 6.64783607365e-12
R_1_115 n679 PAR_2_1_VSS 0.371152097236
L_2_115 PAR_1_2_VDD075CPU n680 3.13090536726e-11
R_2_115 n680 PAR_2_1_VSS 0.370555633404
R_3_115 PAR_1_2_VDD075CPU n681 0.14334240579
C_3_115 n681 PAR_2_1_VSS 7.19066488768e-10
L_4_115 PAR_1_2_VDD075CPU n682 1.75370153527e-09
R_4_115 n682 PAR_2_1_VSS 9.04559611136
L_5_115 PAR_1_2_VDD075CPU n683 4.53745138665e-07
R_5_115 n683 PAR_2_1_VSS 146.587832309
L_6_115 PAR_1_2_VDD075CPU n684 4.21756277361e-06
R_6_115 n684 PAR_2_1_VSS 334.038057697
R0_116 PAR_1_2_VDD075CPU PAR_2_1_VDD075CPU 0.340946711696
C0_116 PAR_1_2_VDD075CPU PAR_2_1_VDD075CPU 1.40365110098e-10
L_1_116 PAR_1_2_VDD075CPU n685 6.27248450309e-12
R_1_116 n685 PAR_2_1_VDD075CPU 0.307438974175
L_2_116 PAR_1_2_VDD075CPU n686 4.13495510295e-11
R_2_116 n686 PAR_2_1_VDD075CPU 0.373059341509
L_3_116 PAR_1_2_VDD075CPU n687 1.83883703961e-08
R_3_116 n687 PAR_2_1_VDD075CPU 46.4123481662
L_4_116 PAR_1_2_VDD075CPU n688 1.94297258587e-07
R_4_116 n688 PAR_2_1_VDD075CPU 186.973371389
L_5_116 PAR_1_2_VDD075CPU n689 5.58056264736e-06
R_5_116 n689 PAR_2_1_VDD075CPU 949.583249268
R_6_116 PAR_1_2_VDD075CPU n690 9286.3307524
C_6_116 n690 PAR_2_1_VDD075CPU 1.52098125976e-10
G0_117 PAR_1_2_VDD075CPU PAR_0_2_VSS PAR_1_2_VDD075CPU PAR_0_2_VSS -0.0677015718821
C0_117 PAR_1_2_VDD075CPU PAR_0_2_VSS 1.81327000523e-10
R_1_117 PAR_1_2_VDD075CPU n691 0.0248556557961
C_1_117 n691 PAR_0_2_VSS 6.21114489926e-10
R_2_117 PAR_1_2_VDD075CPU n692 0.0187975930924
C_2_117 n692 PAR_0_2_VSS 2.00421485561e-09
R_3_117 PAR_1_2_VDD075CPU n693 0.0383984906355
C_3_117 n693 PAR_0_2_VSS 2.61408075301e-09
L_4_117 PAR_1_2_VDD075CPU n694 8.44006807703e-09
R_4_117 n694 PAR_0_2_VSS 14.7707052772
R_5_117 PAR_1_2_VDD075CPU n695 30.5734650872
C_5_117 n695 PAR_0_2_VSS 1.90501784404e-10
R_6_117 PAR_1_2_VDD075CPU n696 91.7223108445
C_6_117 n696 PAR_0_2_VSS 1.79262526117e-10
R0_118 PAR_1_2_VDD075CPU PAR_0_2_VDD075CPU 0.00396624737025
C0_118 PAR_1_2_VDD075CPU PAR_0_2_VDD075CPU 4.85046402829e-11
L_1_118 PAR_1_2_VDD075CPU n697 6.38112046193e-13
R_1_118 n697 PAR_0_2_VDD075CPU 0.0394021112582
L_2_118 PAR_1_2_VDD075CPU n698 1.00659810397e-12
R_2_118 n698 PAR_0_2_VDD075CPU 0.0258157997967
L_3_118 PAR_1_2_VDD075CPU n699 5.40262790444e-12
R_3_118 n699 PAR_0_2_VDD075CPU 0.0524158681228
L_4_118 PAR_1_2_VDD075CPU n700 2.08340241695e-08
R_4_118 n700 PAR_0_2_VDD075CPU 42.6342252671
L_5_118 PAR_1_2_VDD075CPU n701 1.505757339e-06
R_5_118 n701 PAR_0_2_VDD075CPU 471.729770563
G0_119 PAR_1_2_VDD075CPU PAR_1_2_VSS PAR_1_2_VDD075CPU PAR_1_2_VSS -0.0163956497709
C0_119 PAR_1_2_VDD075CPU PAR_1_2_VSS 5.69350118611e-11
R_1_119 PAR_1_2_VDD075CPU n702 0.00175919087879
C_1_119 n702 PAR_1_2_VSS 9.76337018155e-09
R_2_119 PAR_1_2_VDD075CPU n703 0.000804044322002
C_2_119 n703 PAR_1_2_VSS 4.65124133283e-08
R_3_119 PAR_1_2_VDD075CPU n704 0.00375977767407
C_3_119 n704 PAR_1_2_VSS 2.48975486701e-08
R_4_119 PAR_1_2_VDD075CPU n705 0.250583262158
C_4_119 n705 PAR_1_2_VSS 5.59054244184e-10
R_5_119 PAR_1_2_VDD075CPU n706 9.75425023683
C_5_119 n706 PAR_1_2_VSS 7.85689917028e-11
L_6_119 PAR_1_2_VDD075CPU n707 5.14051518838e-07
R_6_119 n707 PAR_1_2_VSS 60.9917813997
G0_120 PAR_1_2_VDD075CPU PAR_0_0_VSS PAR_1_2_VDD075CPU PAR_0_0_VSS -0.401631010361
C0_120 PAR_1_2_VDD075CPU PAR_0_0_VSS 2.45085239798e-10
R_1_120 PAR_1_2_VDD075CPU n708 0.0175327924123
C_1_120 n708 PAR_0_0_VSS 7.70300888219e-10
L_2_120 PAR_1_2_VDD075CPU n709 7.04743750741e-10
R_2_120 n709 PAR_0_0_VSS 2.48984756804
R_3_120 PAR_1_2_VDD075CPU n710 7.62061742853
C_3_120 n710 PAR_0_0_VSS 1.13692044081e-10
R_4_120 PAR_1_2_VDD075CPU n711 62.0529061307
C_4_120 n711 PAR_0_0_VSS 1.25465026775e-10
G0_121 PAR_2_2_VSS PAR_0_0_VDD075CPU PAR_2_2_VSS PAR_0_0_VDD075CPU -0.0243527622441
C0_121 PAR_2_2_VSS PAR_0_0_VDD075CPU 2.79577428879e-11
R_1_121 PAR_2_2_VSS n712 0.131067738483
C_1_121 n712 PAR_0_0_VDD075CPU 1.14006768291e-10
R_2_121 PAR_2_2_VSS n713 1.75176268417
C_2_121 n713 PAR_0_0_VDD075CPU 4.42917436893e-11
L_3_121 PAR_2_2_VSS n714 1.75195945614e-07
R_3_121 n714 PAR_0_0_VDD075CPU 48.4499016949
L_4_121 PAR_2_2_VSS n715 5.27806490746e-06
R_4_121 n715 PAR_0_0_VDD075CPU 269.332134859
G0_122 PAR_2_2_VSS PAR_1_0_VSS PAR_2_2_VSS PAR_1_0_VSS -0.272028155874
C0_122 PAR_2_2_VSS PAR_1_0_VSS 3.28809773802e-11
R_1_122 PAR_2_2_VSS n716 0.294136190479
C_1_122 n716 PAR_1_0_VSS 1.17439644702e-10
R_2_122 PAR_2_2_VSS n717 1.53086869578
C_2_122 n717 PAR_1_0_VSS 8.50261265475e-11
R_3_122 PAR_2_2_VSS n718 0.350894982992
C_3_122 n718 PAR_1_0_VSS 7.20602932483e-10
R_4_122 PAR_2_2_VSS n719 0.484680458036
C_4_122 n719 PAR_1_0_VSS 1.7677879005e-09
L_5_122 PAR_2_2_VSS n720 2.25028844838e-08
R_5_122 n720 PAR_1_0_VSS 5.06970530547
L_6_122 PAR_2_2_VSS n721 1.95335240363e-07
R_6_122 n721 PAR_1_0_VSS 13.3729062158
G0_123 PAR_2_2_VSS PAR_1_0_VDD075CPU PAR_2_2_VSS PAR_1_0_VDD075CPU -0.0273497313864
C0_123 PAR_2_2_VSS PAR_1_0_VDD075CPU 4.06771147408e-11
R_1_123 PAR_2_2_VSS n722 0.176689972624
C_1_123 n722 PAR_1_0_VDD075CPU 9.70847943838e-11
R_2_123 PAR_2_2_VSS n723 1.54402874804
C_2_123 n723 PAR_1_0_VDD075CPU 5.371417171e-11
R_3_123 PAR_2_2_VSS n724 87.9671243179
C_3_123 n724 PAR_1_0_VDD075CPU 7.10251738355e-12
L_4_123 PAR_2_2_VSS n725 1.28714133541e-07
R_4_123 n725 PAR_1_0_VDD075CPU 58.1037958836
L_5_123 PAR_2_2_VSS n726 1.00382304973e-06
R_5_123 n726 PAR_1_0_VDD075CPU 98.6275556185
G0_124 PAR_2_2_VSS PAR_2_0_VSS PAR_2_2_VSS PAR_2_0_VSS -0.384247550171
C0_124 PAR_2_2_VSS PAR_2_0_VSS 5.62249447549e-11
R_1_124 PAR_2_2_VSS n727 0.279149557638
C_1_124 n727 PAR_2_0_VSS 1.14647453619e-10
R_2_124 PAR_2_2_VSS n728 1.77519239291
C_2_124 n728 PAR_2_0_VSS 9.76076356798e-11
R_3_124 PAR_2_2_VSS n729 0.324869792753
C_3_124 n729 PAR_2_0_VSS 2.88441693476e-09
L_4_124 PAR_2_2_VSS n730 1.28213978533e-08
R_4_124 n730 PAR_2_0_VSS 3.48358186244
L_5_124 PAR_2_2_VSS n731 1.40994390076e-07
R_5_124 n731 PAR_2_0_VSS 10.2894620339
G0_125 PAR_2_2_VSS PAR_2_0_VDD075CPU PAR_2_2_VSS PAR_2_0_VDD075CPU -0.0326498361456
C0_125 PAR_2_2_VSS PAR_2_0_VDD075CPU 4.59944673214e-11
R_1_125 PAR_2_2_VSS n732 0.176344415866
C_1_125 n732 PAR_2_0_VDD075CPU 1.06142894304e-10
R_2_125 PAR_2_2_VSS n733 1.57548218813
C_2_125 n733 PAR_2_0_VDD075CPU 5.85191000845e-11
R_3_125 PAR_2_2_VSS n734 13.0371512956
C_3_125 n734 PAR_2_0_VDD075CPU 2.39462809435e-11
L_4_125 PAR_2_2_VSS n735 1.07673011042e-07
R_4_125 n735 PAR_2_0_VDD075CPU 46.9872955903
L_5_125 PAR_2_2_VSS n736 9.22445653985e-07
R_5_125 n736 PAR_2_0_VDD075CPU 87.9701673223
R0_126 PAR_2_2_VSS PAR_0_1_VSS 76523.200227
C0_126 PAR_2_2_VSS PAR_0_1_VSS 2.58878259959e-11
R_1_126 PAR_2_2_VSS n737 0.303037679874
C_1_126 n737 PAR_0_1_VSS 1.43954802993e-10
R_2_126 PAR_2_2_VSS n738 0.438760125206
C_2_126 n738 PAR_0_1_VSS 3.70221481384e-10
R_3_126 PAR_2_2_VSS n739 0.424335969484
C_3_126 n739 PAR_0_1_VSS 8.91808701137e-10
R_4_126 PAR_2_2_VSS n740 0.754004254325
C_4_126 n740 PAR_0_1_VSS 1.30045154417e-09
R_5_126 PAR_2_2_VSS n741 1.44673399631
C_5_126 n741 PAR_0_1_VSS 2.56815897957e-09
R_6_126 PAR_2_2_VSS n742 4.26163170813
C_6_126 n742 PAR_0_1_VSS 3.21551731931e-09
G0_127 PAR_2_2_VSS PAR_0_1_VDD075CPU PAR_2_2_VSS PAR_0_1_VDD075CPU -0.0181385772258
C0_127 PAR_2_2_VSS PAR_0_1_VDD075CPU 3.32746926039e-11
R_1_127 PAR_2_2_VSS n743 0.226025366154
C_1_127 n743 PAR_0_1_VDD075CPU 8.37523029052e-11
R_2_127 PAR_2_2_VSS n744 2.93663053091
C_2_127 n744 PAR_0_1_VDD075CPU 3.1233270925e-11
R_3_127 PAR_2_2_VSS n745 37.6079968445
C_3_127 n745 PAR_0_1_VDD075CPU 1.0069518689e-11
L_4_127 PAR_2_2_VSS n746 2.74563729938e-07
R_4_127 n746 PAR_0_1_VDD075CPU 75.2914301081
L_5_127 PAR_2_2_VSS n747 2.91831234016e-06
R_5_127 n747 PAR_0_1_VDD075CPU 205.894533159
R0_128 PAR_2_2_VSS PAR_1_1_VSS 0.179805582476
C0_128 PAR_2_2_VSS PAR_1_1_VSS 1.79999658431e-11
R_1_128 PAR_2_2_VSS n748 0.253007379358
C_1_128 n748 PAR_1_1_VSS 5.10668849033e-11
R_2_128 PAR_2_2_VSS n749 0.811149310596
C_2_128 n749 PAR_1_1_VSS 1.01773460393e-10
L_3_128 PAR_2_2_VSS n750 3.9551118303e-11
R_3_128 n750 PAR_1_1_VSS 0.364646356034
R_4_128 PAR_2_2_VSS n751 50.229191077
C_4_128 n751 PAR_1_1_VSS 7.31180393005e-12
L_5_128 PAR_2_2_VSS n752 4.38421919645e-07
R_5_128 n752 PAR_1_1_VSS 133.50232667
L_6_128 PAR_2_2_VSS n753 3.64805614686e-06
R_6_128 n753 PAR_1_1_VSS 288.348316927
G0_129 PAR_2_2_VSS PAR_1_1_VDD075CPU PAR_2_2_VSS PAR_1_1_VDD075CPU -0.0124943783976
C0_129 PAR_2_2_VSS PAR_1_1_VDD075CPU 1.68901430704e-11
R_1_129 PAR_2_2_VSS n754 0.190522809848
C_1_129 n754 PAR_1_1_VDD075CPU 6.25721121177e-11
R_2_129 PAR_2_2_VSS n755 0.531325296458
C_2_129 n755 PAR_1_1_VDD075CPU 2.26394063207e-10
R_3_129 PAR_2_2_VSS n756 65.5552539534
C_3_129 n756 PAR_1_1_VDD075CPU 9.55296975661e-12
L_4_129 PAR_2_2_VSS n757 4.53859756329e-07
R_4_129 n757 PAR_1_1_VDD075CPU 80.035979724
R0_130 PAR_2_2_VSS PAR_2_1_VSS 0.021441548448
L_1_130 PAR_2_2_VSS n758 1.69731429884e-11
R_1_130 n758 PAR_2_1_VSS 0.388438893401
L_2_130 PAR_2_2_VSS n759 1.88401680108e-11
R_2_130 n759 PAR_2_1_VSS 0.152459353983
L_3_130 PAR_2_2_VSS n760 4.17520682194e-11
R_3_130 n760 PAR_2_1_VSS 0.141085630515
L_4_130 PAR_2_2_VSS n761 1.95187828985e-10
R_4_130 n761 PAR_2_1_VSS 0.291864115033
L_5_130 PAR_2_2_VSS n762 2.62030630638e-09
R_5_130 n762 PAR_2_1_VSS 1.6156287342
L_6_130 PAR_2_2_VSS n763 1.81354133038e-07
R_6_130 n763 PAR_2_1_VSS 18.8189254552
G0_131 PAR_2_2_VSS PAR_2_1_VDD075CPU PAR_2_2_VSS PAR_2_1_VDD075CPU -0.0096147258011
C0_131 PAR_2_2_VSS PAR_2_1_VDD075CPU 3.23818582305e-11
R_1_131 PAR_2_2_VSS n764 0.224205494698
C_1_131 n764 PAR_2_1_VDD075CPU 8.98675438065e-11
R_2_131 PAR_2_2_VSS n765 0.443572271913
C_2_131 n765 PAR_2_1_VDD075CPU 1.89825413596e-10
R_3_131 PAR_2_2_VSS n766 0.970967398028
C_3_131 n766 PAR_2_1_VDD075CPU 1.94812489779e-10
R_4_131 PAR_2_2_VSS n767 2.69000955929
C_4_131 n767 PAR_2_1_VDD075CPU 1.49480582248e-10
R_5_131 PAR_2_2_VSS n768 17.8673068152
C_5_131 n768 PAR_2_1_VDD075CPU 5.37969957313e-11
L_6_131 PAR_2_2_VSS n769 9.01668134732e-07
R_6_131 n769 PAR_2_1_VDD075CPU 104.007100721
R0_132 PAR_2_2_VSS PAR_0_2_VSS 1637.63584614
C0_132 PAR_2_2_VSS PAR_0_2_VSS 2.59721941112e-11
R_1_132 PAR_2_2_VSS n770 0.339653953731
C_1_132 n770 PAR_0_2_VSS 1.31166667139e-10
R_2_132 PAR_2_2_VSS n771 0.452245033952
C_2_132 n771 PAR_0_2_VSS 3.45969521611e-10
R_3_132 PAR_2_2_VSS n772 0.493508452723
C_3_132 n772 PAR_0_2_VSS 7.74051422197e-10
R_4_132 PAR_2_2_VSS n773 0.753738769522
C_4_132 n773 PAR_0_2_VSS 1.31816544813e-09
R_5_132 PAR_2_2_VSS n774 1.55791798732
C_5_132 n774 PAR_0_2_VSS 2.53400453363e-09
R_6_132 PAR_2_2_VSS n775 4.61319295247
C_6_132 n775 PAR_0_2_VSS 2.93641106558e-09
G0_133 PAR_2_2_VSS PAR_0_2_VDD075CPU PAR_2_2_VSS PAR_0_2_VDD075CPU -0.020847360414
C0_133 PAR_2_2_VSS PAR_0_2_VDD075CPU 3.22596764222e-11
R_1_133 PAR_2_2_VSS n776 0.174419116471
C_1_133 n776 PAR_0_2_VDD075CPU 1.02863845061e-10
R_2_133 PAR_2_2_VSS n777 2.4570039832
C_2_133 n777 PAR_0_2_VDD075CPU 3.11982227146e-11
L_3_133 PAR_2_2_VSS n778 2.18787659015e-07
R_3_133 n778 PAR_0_2_VDD075CPU 75.0502322062
L_4_133 PAR_2_2_VSS n779 1.46420937779e-06
R_4_133 n779 PAR_0_2_VDD075CPU 149.509946184
L_5_133 PAR_2_2_VSS n780 3.04484984482e-05
R_5_133 n780 PAR_0_2_VDD075CPU 1198.4149611
R0_134 PAR_2_2_VSS PAR_1_2_VSS 0.0113566919992
L_1_134 PAR_2_2_VSS n781 3.68004742262e-12
R_1_134 n781 PAR_1_2_VSS 0.079894940087
L_2_134 PAR_2_2_VSS n782 6.95764647654e-12
R_2_134 n782 PAR_1_2_VSS 0.0584451056987
L_3_134 PAR_2_2_VSS n783 1.17182303966e-10
R_3_134 n783 PAR_1_2_VSS 0.305557019094
L_4_134 PAR_2_2_VSS n784 1.51854869825e-10
R_4_134 n784 PAR_1_2_VSS 0.172450855334
L_5_134 PAR_2_2_VSS n785 1.72056609841e-09
R_5_134 n785 PAR_1_2_VSS 0.809238568879
L_6_134 PAR_2_2_VSS n786 9.88001994032e-08
R_6_134 n786 PAR_1_2_VSS 9.38570493023
G0_135 PAR_2_2_VSS PAR_1_2_VDD075CPU PAR_2_2_VSS PAR_1_2_VDD075CPU -0.0143760102761
C0_135 PAR_2_2_VSS PAR_1_2_VDD075CPU 3.32874054238e-11
R_1_135 PAR_2_2_VSS n787 0.184683261728
C_1_135 n787 PAR_1_2_VDD075CPU 1.09392804621e-10
R_2_135 PAR_2_2_VSS n788 0.0434839840413
C_2_135 n788 PAR_1_2_VDD075CPU 2.36222973386e-09
R_3_135 PAR_2_2_VSS n789 3.29436525643
C_3_135 n789 PAR_1_2_VDD075CPU 4.95108437309e-11
R_4_135 PAR_2_2_VSS n790 13.7019122189
C_4_135 n790 PAR_1_2_VDD075CPU 4.37500085697e-11
L_5_135 PAR_2_2_VSS n791 4.67727381389e-07
R_5_135 n791 PAR_1_2_VDD075CPU 94.4136744603
L_6_135 PAR_2_2_VSS n792 4.11225479368e-06
R_6_135 n792 PAR_1_2_VDD075CPU 264.247832956
R0_136 PAR_2_2_VSS PAR_0_0_VSS 164961.356152
R_1_136 PAR_2_2_VSS n793 0.053203181771
C_1_136 n793 PAR_0_0_VSS 6.90058809496e-10
R_2_136 PAR_2_2_VSS n794 0.179829069879
C_2_136 n794 PAR_0_0_VSS 7.51838447182e-10
R_3_136 PAR_2_2_VSS n795 0.29803979651
C_3_136 n795 PAR_0_0_VSS 1.03074889714e-09
R_4_136 PAR_2_2_VSS n796 0.22604714823
C_4_136 n796 PAR_0_0_VSS 4.69085769288e-09
R_5_136 PAR_2_2_VSS n797 0.640251652521
C_5_136 n797 PAR_0_0_VSS 3.79497403165e-09
R_6_136 PAR_2_2_VSS n798 6.56403689415
C_6_136 n798 PAR_0_0_VSS 1.7857314902e-09
G0_137 PAR_2_2_VDD075CPU PAR_0_0_VDD075CPU PAR_2_2_VDD075CPU PAR_0_0_VDD075CPU -0.393018733893
C0_137 PAR_2_2_VDD075CPU PAR_0_0_VDD075CPU 1.96259008371e-11
R_1_137 PAR_2_2_VDD075CPU n799 4.25906143317
C_1_137 n799 PAR_0_0_VDD075CPU 5.95317557489e-12
L_2_137 PAR_2_2_VDD075CPU n800 3.5799726537e-10
R_2_137 n800 PAR_0_0_VDD075CPU 3.32155994314
R_3_137 PAR_2_2_VDD075CPU n801 8.20791691028
C_3_137 n801 PAR_0_0_VDD075CPU 2.62929130061e-11
L_4_137 PAR_2_2_VDD075CPU n802 5.69443529828e-09
R_4_137 n802 PAR_0_0_VDD075CPU 12.4146548725
R_5_137 PAR_2_2_VDD075CPU n803 28.9239399709
C_5_137 n803 PAR_0_0_VDD075CPU 3.62549336772e-11
L_6_137 PAR_2_2_VDD075CPU n804 3.03524296732e-07
R_6_137 n804 PAR_0_0_VDD075CPU 87.803208095
R_7_137 PAR_2_2_VDD075CPU n805 549.997066128
C_7_137 n805 PAR_0_0_VDD075CPU 2.51546822992e-11
G0_138 PAR_2_2_VDD075CPU PAR_1_0_VSS PAR_2_2_VDD075CPU PAR_1_0_VSS -0.125226411476
C0_138 PAR_2_2_VDD075CPU PAR_1_0_VSS 2.20848916907e-11
R_1_138 PAR_2_2_VDD075CPU n806 1.69363354026
C_1_138 n806 PAR_1_0_VSS 1.80058867216e-11
R_2_138 PAR_2_2_VDD075CPU n807 2.37865047239
C_2_138 n807 PAR_1_0_VSS 3.69190126411e-11
L_3_138 PAR_2_2_VDD075CPU n808 2.68012934522e-09
R_3_138 n808 PAR_1_0_VSS 9.55921660136
L_4_138 PAR_2_2_VDD075CPU n809 6.48753570093e-08
R_4_138 n809 PAR_1_0_VSS 54.4925258364
L_5_138 PAR_2_2_VDD075CPU n810 2.81444936574e-06
R_5_138 n810 PAR_1_0_VSS 618.689668282
L_6_138 PAR_2_2_VDD075CPU n811 2.37976150281e-05
R_6_138 n811 PAR_1_0_VSS 1543.51690825
G0_139 PAR_2_2_VDD075CPU PAR_1_0_VDD075CPU PAR_2_2_VDD075CPU PAR_1_0_VDD075CPU -0.171590675443
C0_139 PAR_2_2_VDD075CPU PAR_1_0_VDD075CPU 2.08466795961e-11
R_1_139 PAR_2_2_VDD075CPU n812 5.87968052926
C_1_139 n812 PAR_1_0_VDD075CPU 1.54459937993e-12
L_2_139 PAR_2_2_VDD075CPU n813 6.77230022394e-10
R_2_139 n813 PAR_1_0_VDD075CPU 5.9421003358
R_3_139 PAR_2_2_VDD075CPU n814 876.32245917
C_3_139 n814 PAR_1_0_VDD075CPU 5.16689677625e-13
L_4_139 PAR_2_2_VDD075CPU n815 5.8669971095e-07
R_4_139 n815 PAR_1_0_VDD075CPU 316.070850813
R_5_139 PAR_2_2_VDD075CPU n816 2686.1849946
C_5_139 n816 PAR_1_0_VDD075CPU 5.70285164234e-12
L_6_139 PAR_2_2_VDD075CPU n817 0.259193602994
R_6_139 n817 PAR_1_0_VDD075CPU 6058.67091637
G0_140 PAR_2_2_VDD075CPU PAR_2_0_VSS PAR_2_2_VDD075CPU PAR_2_0_VSS -0.0298621530693
C0_140 PAR_2_2_VDD075CPU PAR_2_0_VSS 2.59941356407e-11
R_1_140 PAR_2_2_VDD075CPU n818 3.91884391791
C_1_140 n818 PAR_2_0_VSS 9.32315128553e-12
R_2_140 PAR_2_2_VDD075CPU n819 9.88365880734
C_2_140 n819 PAR_2_0_VSS 8.28286905101e-12
R_3_140 PAR_2_2_VDD075CPU n820 35.1933165003
C_3_140 n820 PAR_2_0_VSS 1.69889428277e-11
L_4_140 PAR_2_2_VDD075CPU n821 4.39081230584e-08
R_4_140 n821 PAR_2_0_VSS 37.5139187335
L_5_140 PAR_2_2_VDD075CPU n822 1.55559094514e-06
R_5_140 n822 PAR_2_0_VSS 428.272943537
L_6_140 PAR_2_2_VDD075CPU n823 1.63250195644e-05
R_6_140 n823 PAR_2_0_VSS 1148.86634908
G0_141 PAR_2_2_VDD075CPU PAR_2_0_VDD075CPU PAR_2_2_VDD075CPU PAR_2_0_VDD075CPU -0.175721579352
C0_141 PAR_2_2_VDD075CPU PAR_2_0_VDD075CPU 2.24630434806e-11
R_1_141 PAR_2_2_VDD075CPU n824 5.73415400752
C_1_141 n824 PAR_2_0_VDD075CPU 1.88239481299e-12
L_2_141 PAR_2_2_VDD075CPU n825 6.77751775248e-10
R_2_141 n825 PAR_2_0_VDD075CPU 5.87299671159
R_3_141 PAR_2_2_VDD075CPU n826 859.436640459
C_3_141 n826 PAR_2_0_VDD075CPU 4.00121446997e-13
L_4_141 PAR_2_2_VDD075CPU n827 1.76939453786e-07
R_4_141 n827 PAR_2_0_VDD075CPU 183.206177495
R_5_141 PAR_2_2_VDD075CPU n828 6083.29308923
C_5_141 n828 PAR_2_0_VDD075CPU 1.43626541124e-12
G0_142 PAR_2_2_VDD075CPU PAR_0_1_VSS PAR_2_2_VDD075CPU PAR_0_1_VSS -0.113477578097
C0_142 PAR_2_2_VDD075CPU PAR_0_1_VSS 2.1041813023e-11
R_1_142 PAR_2_2_VDD075CPU n829 1.31801007168
C_1_142 n829 PAR_0_1_VSS 1.95694044538e-11
R_2_142 PAR_2_2_VDD075CPU n830 1.41504573476
C_2_142 n830 PAR_0_1_VSS 5.28772291141e-11
L_3_142 PAR_2_2_VDD075CPU n831 2.87884084817e-09
R_3_142 n831 PAR_0_1_VSS 11.2284039105
L_4_142 PAR_2_2_VDD075CPU n832 2.90545886485e-08
R_4_142 n832 PAR_0_1_VSS 40.9538517451
R_5_142 PAR_2_2_VDD075CPU n833 339.068323373
C_5_142 n833 PAR_0_1_VSS 1.76532872774e-11
R_6_142 PAR_2_2_VDD075CPU n834 670.416863319
C_6_142 n834 PAR_0_1_VSS 2.42134163319e-11
G0_143 PAR_2_2_VDD075CPU PAR_0_1_VDD075CPU PAR_2_2_VDD075CPU PAR_0_1_VDD075CPU -0.477544334368
C0_143 PAR_2_2_VDD075CPU PAR_0_1_VDD075CPU 1.43392600108e-11
R_1_143 PAR_2_2_VDD075CPU n835 3.2822105186
C_1_143 n835 PAR_0_1_VDD075CPU 1.46984379874e-11
L_2_143 PAR_2_2_VDD075CPU n836 2.53707555282e-10
R_2_143 n836 PAR_0_1_VDD075CPU 2.4069203999
R_3_143 PAR_2_2_VDD075CPU n837 6.38506142309
C_3_143 n837 PAR_0_1_VDD075CPU 3.25872860301e-11
L_4_143 PAR_2_2_VDD075CPU n838 9.7060815281e-09
R_4_143 n838 PAR_0_1_VDD075CPU 17.4190323
R_5_143 PAR_2_2_VDD075CPU n839 61.5155525467
C_5_143 n839 PAR_0_1_VDD075CPU 3.23011731726e-11
L_6_143 PAR_2_2_VDD075CPU n840 2.50683866648e-06
R_6_143 n840 PAR_0_1_VDD075CPU 214.494674554
G0_144 PAR_2_2_VDD075CPU PAR_1_1_VSS PAR_2_2_VDD075CPU PAR_1_1_VSS -0.618981876797
C0_144 PAR_2_2_VDD075CPU PAR_1_1_VSS 1.16912242338e-11
L_1_144 PAR_2_2_VDD075CPU n841 1.25557949096e-10
R_1_144 n841 PAR_1_1_VSS 1.70156883518
R_2_144 PAR_2_2_VDD075CPU n842 0.380106893165
C_2_144 n842 PAR_1_1_VSS 2.93270676698e-10
L_3_144 PAR_2_2_VDD075CPU n843 6.62616862578e-09
R_3_144 n843 PAR_1_1_VSS 32.3625733166
L_4_144 PAR_2_2_VDD075CPU n844 5.00725058434e-06
R_4_144 n844 PAR_1_1_VSS 2570.41327893
R0_145 PAR_2_2_VDD075CPU PAR_1_1_VDD075CPU 0.175124347376
C0_145 PAR_2_2_VDD075CPU PAR_1_1_VDD075CPU 9.61298283135e-12
L_1_145 PAR_2_2_VDD075CPU n845 6.8868614251e-11
R_1_145 n845 PAR_1_1_VDD075CPU 2.90344944373
R_2_145 PAR_2_2_VDD075CPU n846 1.15360942195
C_2_145 n846 PAR_1_1_VDD075CPU 7.15709046782e-11
L_3_145 PAR_2_2_VDD075CPU n847 3.27440414637e-11
R_3_145 n847 PAR_1_1_VDD075CPU 0.305007035559
L_4_145 PAR_2_2_VDD075CPU n848 4.04139026889e-07
R_4_145 n848 PAR_1_1_VDD075CPU 569.991785483
G0_146 PAR_2_2_VDD075CPU PAR_2_1_VSS PAR_2_2_VDD075CPU PAR_2_1_VSS -0.000486248042813
C0_146 PAR_2_2_VDD075CPU PAR_2_1_VSS 2.34055423277e-11
R_1_146 PAR_2_2_VDD075CPU n849 0.17438020785
C_1_146 n849 PAR_2_1_VSS 7.11685562993e-11
R_2_146 PAR_2_2_VDD075CPU n850 0.507146311272
C_2_146 n850 PAR_2_1_VSS 1.23526363703e-10
R_3_146 PAR_2_2_VDD075CPU n851 0.137566351159
C_3_146 n851 PAR_2_1_VSS 7.29377332432e-10
R_4_146 PAR_2_2_VDD075CPU n852 9.11338271237
C_4_146 n852 PAR_2_1_VSS 3.54740163199e-11
R_5_146 PAR_2_2_VDD075CPU n853 39.1631454835
C_5_146 n853 PAR_2_1_VSS 1.89826006679e-11
L_6_146 PAR_2_2_VDD075CPU n854 2.09516201607e-05
R_6_146 n854 PAR_2_1_VSS 2056.55369297
R0_147 PAR_2_2_VDD075CPU PAR_2_1_VDD075CPU 0.0268064312373
L_1_147 PAR_2_2_VDD075CPU n855 2.74724173306e-12
R_1_147 n855 PAR_2_1_VDD075CPU 0.210350012334
L_2_147 PAR_2_2_VDD075CPU n856 7.1903708519e-11
R_2_147 n856 PAR_2_1_VDD075CPU 1.13075991219
L_3_147 PAR_2_2_VDD075CPU n857 2.31681953801e-11
R_3_147 n857 PAR_2_1_VDD075CPU 0.232757560821
R_4_147 PAR_2_2_VDD075CPU n858 647.815671653
C_4_147 n858 PAR_2_1_VDD075CPU 5.16729636772e-13
L_5_147 PAR_2_2_VDD075CPU n859 2.60633741744e-07
R_5_147 n859 PAR_2_1_VDD075CPU 210.668788417
R_6_147 PAR_2_2_VDD075CPU n860 1218.12396915
C_6_147 n860 PAR_2_1_VDD075CPU 3.24545627579e-11
G0_148 PAR_2_2_VDD075CPU PAR_0_2_VSS PAR_2_2_VDD075CPU PAR_0_2_VSS -0.108766168296
C0_148 PAR_2_2_VDD075CPU PAR_0_2_VSS 1.97677209004e-11
R_1_148 PAR_2_2_VDD075CPU n861 1.52938627637
C_1_148 n861 PAR_0_2_VSS 1.5940835728e-11
R_2_148 PAR_2_2_VDD075CPU n862 1.41910510851
C_2_148 n862 PAR_0_2_VSS 5.08974748364e-11
L_3_148 PAR_2_2_VDD075CPU n863 2.73055456126e-09
R_3_148 n863 PAR_0_2_VSS 11.4043935572
L_4_148 PAR_2_2_VDD075CPU n864 3.46350468357e-08
R_4_148 n864 PAR_0_2_VSS 47.4368300507
R_5_148 PAR_2_2_VDD075CPU n865 310.890315135
C_5_148 n865 PAR_0_2_VSS 2.09317344101e-11
R_6_148 PAR_2_2_VDD075CPU n866 910.542750141
C_6_148 n866 PAR_0_2_VSS 1.90823883542e-11
G0_149 PAR_2_2_VDD075CPU PAR_0_2_VDD075CPU PAR_2_2_VDD075CPU PAR_0_2_VDD075CPU -0.184010154504
C0_149 PAR_2_2_VDD075CPU PAR_0_2_VDD075CPU 1.97594232078e-11
R_1_149 PAR_2_2_VDD075CPU n867 5.29313681096
C_1_149 n867 PAR_0_2_VDD075CPU 1.52077818106e-12
L_2_149 PAR_2_2_VDD075CPU n868 7.2094875383e-10
R_2_149 n868 PAR_0_2_VDD075CPU 8.43588348373
L_3_149 PAR_2_2_VDD075CPU n869 2.05045677271e-09
R_3_149 n869 PAR_0_2_VDD075CPU 16.0137731738
L_4_149 PAR_2_2_VDD075CPU n870 1.74163776718e-07
R_4_149 n870 PAR_0_2_VDD075CPU 370.132862597
L_5_149 PAR_2_2_VDD075CPU n871 3.8147491494e-06
R_5_149 n871 PAR_0_2_VDD075CPU 2165.91753138
G0_150 PAR_2_2_VDD075CPU PAR_1_2_VSS PAR_2_2_VDD075CPU PAR_1_2_VSS -2.14725097236
C0_150 PAR_2_2_VDD075CPU PAR_1_2_VSS 1.6005835216e-11
L_1_150 PAR_2_2_VDD075CPU n872 2.6443527185e-11
R_1_150 n872 PAR_1_2_VSS 0.46595559678
R_2_150 PAR_2_2_VDD075CPU n873 0.0794972534429
C_2_150 n873 PAR_1_2_VSS 1.33003810838e-09
R_3_150 PAR_2_2_VDD075CPU n874 3.95016292447
C_3_150 n874 PAR_1_2_VSS 5.55057685367e-11
R_4_150 PAR_2_2_VDD075CPU n875 15.8969933569
C_4_150 n875 PAR_1_2_VSS 5.25117582553e-11
L_5_150 PAR_2_2_VDD075CPU n876 1.12878914611e-05
R_5_150 n876 PAR_1_2_VSS 889.891899047
R0_151 PAR_2_2_VDD075CPU PAR_1_2_VDD075CPU 0.0095842890722
C0_151 PAR_2_2_VDD075CPU PAR_1_2_VDD075CPU 3.2425852145e-11
L_1_151 PAR_2_2_VDD075CPU n877 1.84233533763e-12
R_1_151 n877 PAR_1_2_VDD075CPU 0.108026030297
L_2_151 PAR_2_2_VDD075CPU n878 6.28095878395e-12
R_2_151 n878 PAR_1_2_VDD075CPU 0.0569943671008
R_3_151 PAR_2_2_VDD075CPU n879 3.57317574269
C_3_151 n879 PAR_1_2_VDD075CPU 1.31897486997e-10
L_4_151 PAR_2_2_VDD075CPU n880 9.83249799264e-08
R_4_151 n880 PAR_1_2_VDD075CPU 22.749449362
R_1_152 PAR_2_2_VDD075CPU n881 0.158836135071
C_1_152 n881 PAR_2_2_VSS 5.15204254742e-11
R_2_152 PAR_2_2_VDD075CPU n882 0.0584928600919
C_2_152 n882 PAR_2_2_VSS 1.32711930128e-09
R_3_152 PAR_2_2_VDD075CPU n883 0.0170250220461
C_3_152 n883 PAR_2_2_VSS 5.83468479743e-09
R_4_152 PAR_2_2_VDD075CPU n884 4.29148673618
C_4_152 n884 PAR_2_2_VSS 7.68646097994e-11
R_5_152 PAR_2_2_VDD075CPU n885 29.5910691639
C_5_152 n885 PAR_2_2_VSS 2.70535162288e-11
R_6_152 PAR_2_2_VDD075CPU n886 373.46908563
C_6_152 n886 PAR_2_2_VSS 2.8314631054e-11
G0_153 PAR_2_2_VDD075CPU PAR_0_0_VSS PAR_2_2_VDD075CPU PAR_0_0_VSS -0.304784840094
C0_153 PAR_2_2_VDD075CPU PAR_0_0_VSS 2.64343455892e-11
R_1_153 PAR_2_2_VDD075CPU n887 0.168141845089
C_1_153 n887 PAR_0_0_VSS 9.63547008136e-11
R_2_153 PAR_2_2_VDD075CPU n888 0.599468999155
C_2_153 n888 PAR_0_0_VSS 8.58101825329e-11
L_3_153 PAR_2_2_VDD075CPU n889 7.62037341386e-10
R_3_153 n889 PAR_0_0_VSS 3.48110983644
L_4_153 PAR_2_2_VDD075CPU n890 5.64630522787e-08
R_4_153 n890 PAR_0_0_VSS 57.0771865307
R_5_153 PAR_2_2_VDD075CPU n891 1738.83687256
C_5_153 n891 PAR_0_0_VSS 1.08039378357e-11
G0_154 PAR_0_3_VSS PAR_0_0_VDD075CPU PAR_0_3_VSS PAR_0_0_VDD075CPU -0.199878523726
C0_154 PAR_0_3_VSS PAR_0_0_VDD075CPU 2.01689466742e-10
R_1_154 PAR_0_3_VSS n892 0.0671589059373
C_1_154 n892 PAR_0_0_VDD075CPU 2.67538644294e-10
R_2_154 PAR_0_3_VSS n893 0.220889476208
C_2_154 n893 PAR_0_0_VDD075CPU 3.36671871169e-10
R_3_154 PAR_0_3_VSS n894 1.48502648078
C_3_154 n894 PAR_0_0_VDD075CPU 9.44768888656e-11
L_4_154 PAR_0_3_VSS n895 4.02886665757e-09
R_4_154 n895 PAR_0_0_VDD075CPU 5.00303868592
R_5_154 PAR_0_3_VSS n896 26.8094441564
C_5_154 n896 PAR_0_0_VDD075CPU 2.53296946231e-10
R_6_154 PAR_0_3_VSS n897 132.206932735
C_6_154 n897 PAR_0_0_VDD075CPU 1.49804754302e-10
R0_155 PAR_0_3_VSS PAR_1_0_VSS 70.3421394369
C0_155 PAR_0_3_VSS PAR_1_0_VSS 2.02196620549e-10
R_1_155 PAR_0_3_VSS n898 0.269497160336
C_1_155 n898 PAR_1_0_VSS 1.51457279093e-10
R_2_155 PAR_0_3_VSS n899 0.121500341626
C_2_155 n899 PAR_1_0_VSS 1.79033026857e-09
R_3_155 PAR_0_3_VSS n900 0.104672099491
C_3_155 n900 PAR_1_0_VSS 2.89291187212e-09
R_4_155 PAR_0_3_VSS n901 0.157750930777
C_4_155 n901 PAR_1_0_VSS 4.86187871005e-09
R_5_155 PAR_0_3_VSS n902 1.48576906688
C_5_155 n902 PAR_1_0_VSS 3.5018825887e-09
R_6_155 PAR_0_3_VSS n903 3.76421365499
C_6_155 n903 PAR_1_0_VSS 3.97651635482e-09
G0_156 PAR_0_3_VSS PAR_1_0_VDD075CPU PAR_0_3_VSS PAR_1_0_VDD075CPU -0.196511145976
C0_156 PAR_0_3_VSS PAR_1_0_VDD075CPU 2.31704274723e-10
R_1_156 PAR_0_3_VSS n904 0.0942415837456
C_1_156 n904 PAR_1_0_VDD075CPU 2.11344805328e-10
R_2_156 PAR_0_3_VSS n905 0.210890123734
C_2_156 n905 PAR_1_0_VDD075CPU 3.5438417143e-10
R_3_156 PAR_0_3_VSS n906 1.07003388339
C_3_156 n906 PAR_1_0_VDD075CPU 1.35217239715e-10
L_4_156 PAR_0_3_VSS n907 4.11421155724e-09
R_4_156 n907 PAR_1_0_VDD075CPU 5.08876980528
R_5_156 PAR_0_3_VSS n908 25.2123217117
C_5_156 n908 PAR_1_0_VDD075CPU 2.14178601925e-10
R_6_156 PAR_0_3_VSS n909 59.7530112954
C_6_156 n909 PAR_1_0_VDD075CPU 2.52008060306e-10
R0_157 PAR_0_3_VSS PAR_2_0_VSS 4067.51100724
C0_157 PAR_0_3_VSS PAR_2_0_VSS 2.56581815791e-10
R_1_157 PAR_0_3_VSS n910 0.149837938225
C_1_157 n910 PAR_2_0_VSS 1.68367962099e-10
R_2_157 PAR_0_3_VSS n911 0.342211631876
C_2_157 n911 PAR_2_0_VSS 2.21638363621e-10
R_3_157 PAR_0_3_VSS n912 0.438509417303
C_3_157 n912 PAR_2_0_VSS 6.55744349066e-10
R_4_157 PAR_0_3_VSS n913 0.086141392369
C_4_157 n913 PAR_2_0_VSS 9.3477041032e-09
R_5_157 PAR_0_3_VSS n914 1.40288010518
C_5_157 n914 PAR_2_0_VSS 4.01608713309e-09
R_6_157 PAR_0_3_VSS n915 4.2408298175
C_6_157 n915 PAR_2_0_VSS 3.70251404639e-09
G0_158 PAR_0_3_VSS PAR_2_0_VDD075CPU PAR_0_3_VSS PAR_2_0_VDD075CPU -0.27624846132
C0_158 PAR_0_3_VSS PAR_2_0_VDD075CPU 2.62336148505e-10
R_1_158 PAR_0_3_VSS n916 0.096726153372
C_1_158 n916 PAR_2_0_VDD075CPU 2.6591499348e-10
R_2_158 PAR_0_3_VSS n917 0.216442722877
C_2_158 n917 PAR_2_0_VDD075CPU 4.16065461021e-10
R_3_158 PAR_0_3_VSS n918 1.29605446319
C_3_158 n918 PAR_2_0_VDD075CPU 1.87605324075e-10
L_4_158 PAR_0_3_VSS n919 2.72311059839e-09
R_4_158 n919 PAR_2_0_VDD075CPU 3.61992962902
R_5_158 PAR_0_3_VSS n920 17.1672315279
C_5_158 n920 PAR_2_0_VDD075CPU 4.92059854485e-10
R0_159 PAR_0_3_VSS PAR_0_1_VSS 0.213371965059
C0_159 PAR_0_3_VSS PAR_0_1_VSS 1.7670094253e-10
R_1_159 PAR_0_3_VSS n921 0.337362158221
C_1_159 n921 PAR_0_1_VSS 2.56357094662e-10
R_2_159 PAR_0_3_VSS n922 0.108504833173
C_2_159 n922 PAR_0_1_VSS 1.76456260153e-09
R_3_159 PAR_0_3_VSS n923 0.0752898635516
C_3_159 n923 PAR_0_1_VSS 5.08496481332e-09
R_4_159 PAR_0_3_VSS n924 0.296624502662
C_4_159 n924 PAR_0_1_VSS 2.72974369185e-09
R_5_159 PAR_0_3_VSS n925 0.90010310985
C_5_159 n925 PAR_0_1_VSS 3.41120757497e-09
R_6_159 PAR_0_3_VSS n926 3.98384544283
C_6_159 n926 PAR_0_1_VSS 4.37766875975e-09
G0_160 PAR_0_3_VSS PAR_0_1_VDD075CPU PAR_0_3_VSS PAR_0_1_VDD075CPU -0.1715634902
C0_160 PAR_0_3_VSS PAR_0_1_VDD075CPU 1.92138300576e-10
R_1_160 PAR_0_3_VSS n927 0.118914316434
C_1_160 n927 PAR_0_1_VDD075CPU 2.20765476314e-10
R_2_160 PAR_0_3_VSS n928 0.338390138016
C_2_160 n928 PAR_0_1_VDD075CPU 2.5958271439e-10
R_3_160 PAR_0_3_VSS n929 2.70240590287
C_3_160 n929 PAR_0_1_VDD075CPU 9.01513784001e-11
L_4_160 PAR_0_3_VSS n930 3.94626961235e-09
R_4_160 n930 PAR_0_1_VDD075CPU 5.82874586553
R_5_160 PAR_0_3_VSS n931 25.1406769982
C_5_160 n931 PAR_0_1_VDD075CPU 3.40357738927e-10
G0_161 PAR_0_3_VSS PAR_1_1_VSS PAR_0_3_VSS PAR_1_1_VSS -0.0902770958577
C0_161 PAR_0_3_VSS PAR_1_1_VSS 1.58692086843e-10
R_1_161 PAR_0_3_VSS n932 0.192219803758
C_1_161 n932 PAR_1_1_VSS 1.32265674647e-10
R_2_161 PAR_0_3_VSS n933 1.09488529473
C_2_161 n933 PAR_1_1_VSS 7.47640209712e-11
R_3_161 PAR_0_3_VSS n934 3.93116165295
C_3_161 n934 PAR_1_1_VSS 7.16818141318e-11
L_4_161 PAR_0_3_VSS n935 7.2138612034e-09
R_4_161 n935 PAR_1_1_VSS 11.076632192
R_5_161 PAR_0_3_VSS n936 41.1132757118
C_5_161 n936 PAR_1_1_VSS 2.05422811527e-10
G0_162 PAR_0_3_VSS PAR_1_1_VDD075CPU PAR_0_3_VSS PAR_1_1_VDD075CPU -0.100823366915
C0_162 PAR_0_3_VSS PAR_1_1_VDD075CPU 1.66418213361e-10
R_1_162 PAR_0_3_VSS n937 0.175646786014
C_1_162 n937 PAR_1_1_VDD075CPU 1.49836824021e-10
R_2_162 PAR_0_3_VSS n938 0.635775688644
C_2_162 n938 PAR_1_1_VDD075CPU 1.36472926135e-10
R_3_162 PAR_0_3_VSS n939 2.7774831799
C_3_162 n939 PAR_1_1_VDD075CPU 9.30180239583e-11
L_4_162 PAR_0_3_VSS n940 6.90534961936e-09
R_4_162 n940 PAR_1_1_VDD075CPU 9.91833544645
R_5_162 PAR_0_3_VSS n941 32.7487351517
C_5_162 n941 PAR_1_1_VDD075CPU 2.57342942699e-10
R0_163 PAR_0_3_VSS PAR_2_1_VSS 429.903104164
C0_163 PAR_0_3_VSS PAR_2_1_VSS 2.01926649209e-10
R_1_163 PAR_0_3_VSS n942 0.157782249358
C_1_163 n942 PAR_2_1_VSS 1.83141755808e-10
R_2_163 PAR_0_3_VSS n943 0.510085280302
C_2_163 n943 PAR_2_1_VSS 3.80583894879e-10
R_3_163 PAR_0_3_VSS n944 0.335933698233
C_3_163 n944 PAR_2_1_VSS 1.19419002476e-09
R_4_163 PAR_0_3_VSS n945 1.13737466028
C_4_163 n945 PAR_2_1_VSS 8.8673090171e-10
R_5_163 PAR_0_3_VSS n946 3.07531649632
C_5_163 n946 PAR_2_1_VSS 1.28870945801e-09
R_6_163 PAR_0_3_VSS n947 8.5470317301
C_6_163 n947 PAR_2_1_VSS 1.54243529413e-09
G0_164 PAR_0_3_VSS PAR_2_1_VDD075CPU PAR_0_3_VSS PAR_2_1_VDD075CPU -0.172313883195
C0_164 PAR_0_3_VSS PAR_2_1_VDD075CPU 1.70309572723e-10
R_1_164 PAR_0_3_VSS n948 0.125660591744
C_1_164 n948 PAR_2_1_VDD075CPU 1.62911418982e-10
R_2_164 PAR_0_3_VSS n949 0.299036660392
C_2_164 n949 PAR_2_1_VDD075CPU 2.64690459376e-10
R_3_164 PAR_0_3_VSS n950 1.00780742565
C_3_164 n950 PAR_2_1_VDD075CPU 1.34569852409e-10
L_4_164 PAR_0_3_VSS n951 4.38523724697e-09
R_4_164 n951 PAR_2_1_VDD075CPU 5.80336282715
R_5_164 PAR_0_3_VSS n952 31.3193358289
C_5_164 n952 PAR_2_1_VDD075CPU 2.11551380991e-10
R_6_164 PAR_0_3_VSS n953 138.885790959
C_6_164 n953 PAR_2_1_VDD075CPU 1.37186166369e-10
R0_165 PAR_0_3_VSS PAR_0_2_VSS 0.00640112886876
C0_165 PAR_0_3_VSS PAR_0_2_VSS 1.1498168509e-10
L_1_165 PAR_0_3_VSS n954 4.47950918137e-13
R_1_165 n954 PAR_0_2_VSS 0.0128140443343
R_2_165 PAR_0_3_VSS n955 0.115143522448
C_2_165 n955 PAR_0_2_VSS 2.28247327478e-09
L_3_165 PAR_0_3_VSS n956 1.14860658021e-09
R_3_165 n956 PAR_0_2_VSS 0.393953801236
L_4_165 PAR_0_3_VSS n957 3.70056668924e-09
R_4_165 n957 PAR_0_2_VSS 0.353936664815
G0_166 PAR_0_3_VSS PAR_0_2_VDD075CPU PAR_0_3_VSS PAR_0_2_VDD075CPU -0.0976122232978
C0_166 PAR_0_3_VSS PAR_0_2_VDD075CPU 2.45572499453e-10
R_1_166 PAR_0_3_VSS n958 0.00848270517595
C_1_166 n958 PAR_0_2_VDD075CPU 3.27109135324e-09
R_2_166 PAR_0_3_VSS n959 0.0279316528516
C_2_166 n959 PAR_0_2_VDD075CPU 1.78291393639e-09
R_3_166 PAR_0_3_VSS n960 0.650347072917
C_3_166 n960 PAR_0_2_VDD075CPU 2.56646412724e-10
L_4_166 PAR_0_3_VSS n961 8.11589124065e-09
R_4_166 n961 PAR_0_2_VDD075CPU 10.2446183206
R_5_166 PAR_0_3_VSS n962 20.9626202203
C_5_166 n962 PAR_0_2_VDD075CPU 3.71395028711e-10
R0_167 PAR_0_3_VSS PAR_1_2_VSS 0.127488330877
C0_167 PAR_0_3_VSS PAR_1_2_VSS 1.78373838123e-10
R_1_167 PAR_0_3_VSS n963 0.238323108782
C_1_167 n963 PAR_1_2_VSS 3.55623380835e-10
R_2_167 PAR_0_3_VSS n964 0.218301067563
C_2_167 n964 PAR_1_2_VSS 1.03219395947e-09
R_3_167 PAR_0_3_VSS n965 0.293137481185
C_3_167 n965 PAR_1_2_VSS 2.12149284486e-09
R_4_167 PAR_0_3_VSS n966 0.389766244225
C_4_167 n966 PAR_1_2_VSS 3.58346741305e-09
R_5_167 PAR_0_3_VSS n967 0.95831677377
C_5_167 n967 PAR_1_2_VSS 4.61024294798e-09
R_6_167 PAR_0_3_VSS n968 3.42303381672
C_6_167 n968 PAR_1_2_VSS 4.13045862654e-09
G0_168 PAR_0_3_VSS PAR_1_2_VDD075CPU PAR_0_3_VSS PAR_1_2_VDD075CPU -0.140334004081
C0_168 PAR_0_3_VSS PAR_1_2_VDD075CPU 2.24886603014e-10
R_1_168 PAR_0_3_VSS n969 0.0613900280729
C_1_168 n969 PAR_1_2_VDD075CPU 4.5342602221e-10
R_2_168 PAR_0_3_VSS n970 0.326908319296
C_2_168 n970 PAR_1_2_VDD075CPU 2.37052090454e-10
R_3_168 PAR_0_3_VSS n971 1.86310381929
C_3_168 n971 PAR_1_2_VDD075CPU 1.21692760143e-10
L_4_168 PAR_0_3_VSS n972 5.48454946445e-09
R_4_168 n972 PAR_1_2_VDD075CPU 7.12585656098
R_5_168 PAR_0_3_VSS n973 23.8716507427
C_5_168 n973 PAR_1_2_VDD075CPU 3.5594094029e-10
R0_169 PAR_0_3_VSS PAR_2_2_VSS 128.207722433
C0_169 PAR_0_3_VSS PAR_2_2_VSS 1.60650550955e-11
R_1_169 PAR_0_3_VSS n974 0.275035048219
C_1_169 n974 PAR_2_2_VSS 2.04605740928e-10
R_2_169 PAR_0_3_VSS n975 0.396164056178
C_2_169 n975 PAR_2_2_VSS 4.71261435954e-10
R_3_169 PAR_0_3_VSS n976 0.215490358528
C_3_169 n976 PAR_2_2_VSS 2.13290984729e-09
R_4_169 PAR_0_3_VSS n977 0.456815863385
C_4_169 n977 PAR_2_2_VSS 2.45129809973e-09
R_5_169 PAR_0_3_VSS n978 1.36509793971
C_5_169 n978 PAR_2_2_VSS 2.93934139823e-09
R_6_169 PAR_0_3_VSS n979 4.30351281015
C_6_169 n979 PAR_2_2_VSS 3.09548910794e-09
G0_170 PAR_0_3_VSS PAR_2_2_VDD075CPU PAR_0_3_VSS PAR_2_2_VDD075CPU -0.0869787853211
C0_170 PAR_0_3_VSS PAR_2_2_VDD075CPU 2.36120576341e-11
R_1_170 PAR_0_3_VSS n980 0.973429314777
C_1_170 n980 PAR_2_2_VDD075CPU 2.81779736313e-11
R_2_170 PAR_0_3_VSS n981 0.886534619049
C_2_170 n981 PAR_2_2_VDD075CPU 8.53952909249e-11
L_3_170 PAR_0_3_VSS n982 8.00809587564e-09
R_3_170 n982 PAR_2_2_VDD075CPU 19.6913059811
L_4_170 PAR_0_3_VSS n983 2.35141321989e-08
R_4_170 n983 PAR_2_2_VDD075CPU 27.628160119
R_5_170 PAR_0_3_VSS n984 244.68537144
C_5_170 n984 PAR_2_2_VDD075CPU 3.86973049874e-11
R0_171 PAR_0_3_VSS PAR_0_0_VSS 0.292327359511
C0_171 PAR_0_3_VSS PAR_0_0_VSS 1.54407474726e-10
R_1_171 PAR_0_3_VSS n985 0.0232785987884
C_1_171 n985 PAR_0_0_VSS 1.9089989039e-09
R_2_171 PAR_0_3_VSS n986 0.0426045699828
C_2_171 n986 PAR_0_0_VSS 3.25604907913e-09
R_3_171 PAR_0_3_VSS n987 0.0400096202864
C_3_171 n987 PAR_0_0_VSS 8.37420246934e-09
R_4_171 PAR_0_3_VSS n988 0.0775197343627
C_4_171 n988 PAR_0_0_VSS 1.36024207447e-08
R_5_171 PAR_0_3_VSS n989 0.217993620129
C_5_171 n989 PAR_0_0_VSS 1.97043912134e-08
R_6_171 PAR_0_3_VSS n990 0.282935858753
C_6_171 n990 PAR_0_0_VSS 5.33033787171e-08
G0_172 PAR_0_3_VDD075CPU PAR_0_0_VDD075CPU PAR_0_3_VDD075CPU PAR_0_0_VDD075CPU -10.131691707
C0_172 PAR_0_3_VDD075CPU PAR_0_0_VDD075CPU 1.31876374946e-10
R_1_172 PAR_0_3_VDD075CPU n991 0.317149103881
C_1_172 n991 PAR_0_0_VDD075CPU 1.31244631639e-10
L_2_172 PAR_0_3_VDD075CPU n992 1.34079268755e-11
R_2_172 n992 PAR_0_0_VDD075CPU 0.118190454289
R_3_172 PAR_0_3_VDD075CPU n993 0.157073975326
C_3_172 n993 PAR_0_0_VDD075CPU 9.97172097615e-10
L_4_172 PAR_0_3_VDD075CPU n994 2.74848503889e-10
R_4_172 n994 PAR_0_0_VDD075CPU 0.692027334625
R_5_172 PAR_0_3_VDD075CPU n995 1.75014149014
C_5_172 n995 PAR_0_0_VDD075CPU 6.13655321373e-10
L_6_172 PAR_0_3_VDD075CPU n996 1.57807599014e-08
R_6_172 n996 PAR_0_0_VDD075CPU 4.43326134778
R_7_172 PAR_0_3_VDD075CPU n997 24.5150494667
C_7_172 n997 PAR_0_0_VDD075CPU 5.58043571434e-10
G0_173 PAR_0_3_VDD075CPU PAR_1_0_VSS PAR_0_3_VDD075CPU PAR_1_0_VSS -1.00982518971
C0_173 PAR_0_3_VDD075CPU PAR_1_0_VSS 1.69188594697e-10
R_1_173 PAR_0_3_VDD075CPU n998 0.158924650215
C_1_173 n998 PAR_1_0_VSS 1.67262615075e-10
R_2_173 PAR_0_3_VDD075CPU n999 0.555595837908
C_2_173 n999 PAR_1_0_VSS 2.13855596501e-10
L_3_173 PAR_0_3_VDD075CPU n1000 3.18484991794e-10
R_3_173 n1000 PAR_1_0_VSS 1.10782080444
L_4_173 PAR_0_3_VDD075CPU n1001 1.36945412042e-08
R_4_173 n1001 PAR_1_0_VSS 10.5905603693
L_5_173 PAR_0_3_VDD075CPU n1002 6.51339693371e-07
R_5_173 n1002 PAR_1_0_VSS 78.5643576184
G0_174 PAR_0_3_VDD075CPU PAR_1_0_VDD075CPU PAR_0_3_VDD075CPU PAR_1_0_VDD075CPU -6.05226690164
C0_174 PAR_0_3_VDD075CPU PAR_1_0_VDD075CPU 1.39814609888e-10
R_1_174 PAR_0_3_VDD075CPU n1003 0.215600952385
C_1_174 n1003 PAR_1_0_VDD075CPU 1.77244210097e-10
L_2_174 PAR_0_3_VDD075CPU n1004 1.25374897452e-11
R_2_174 n1004 PAR_1_0_VDD075CPU 0.187394193687
R_3_174 PAR_0_3_VDD075CPU n1005 0.891148777651
C_3_174 n1005 PAR_1_0_VDD075CPU 1.55516753931e-10
L_4_174 PAR_0_3_VDD075CPU n1006 6.0387024333e-10
R_4_174 n1006 PAR_1_0_VDD075CPU 1.64040400974
R_5_174 PAR_0_3_VDD075CPU n1007 3.63796354318
C_5_174 n1007 PAR_1_0_VDD075CPU 2.56935756034e-10
L_6_174 PAR_0_3_VDD075CPU n1008 2.98030964108e-08
R_6_174 n1008 PAR_1_0_VDD075CPU 9.38931920066
R_7_174 PAR_0_3_VDD075CPU n1009 58.6774411735
C_7_174 n1009 PAR_1_0_VDD075CPU 2.22115700818e-10
G0_175 PAR_0_3_VDD075CPU PAR_2_0_VSS PAR_0_3_VDD075CPU PAR_2_0_VSS -0.0913724532617
C0_175 PAR_0_3_VDD075CPU PAR_2_0_VSS 2.01037994795e-10
R_1_175 PAR_0_3_VDD075CPU n1010 0.406708178189
C_1_175 n1010 PAR_2_0_VSS 5.57675036412e-11
R_2_175 PAR_0_3_VDD075CPU n1011 2.70613914297
C_2_175 n1011 PAR_2_0_VSS 5.50590391237e-11
L_3_175 PAR_0_3_VDD075CPU n1012 2.33051439763e-08
R_3_175 n1012 PAR_2_0_VSS 11.4950129468
L_4_175 PAR_0_3_VDD075CPU n1013 5.76843422898e-06
R_4_175 n1013 PAR_2_0_VSS 228.40392684
G0_176 PAR_0_3_VDD075CPU PAR_2_0_VDD075CPU PAR_0_3_VDD075CPU PAR_2_0_VDD075CPU -6.76974087376
C0_176 PAR_0_3_VDD075CPU PAR_2_0_VDD075CPU 1.36465221822e-10
R_1_176 PAR_0_3_VDD075CPU n1014 0.377572458743
C_1_176 n1014 PAR_2_0_VDD075CPU 1.23099854251e-10
L_2_176 PAR_0_3_VDD075CPU n1015 2.40839154651e-11
R_2_176 n1015 PAR_2_0_VDD075CPU 0.18521039594
R_3_176 PAR_0_3_VDD075CPU n1016 0.262574795183
C_3_176 n1016 PAR_2_0_VDD075CPU 8.27971055054e-10
L_4_176 PAR_0_3_VDD075CPU n1017 3.95636281977e-10
R_4_176 n1017 PAR_2_0_VDD075CPU 0.787885729645
R_5_176 PAR_0_3_VDD075CPU n1018 3.2610416216
C_5_176 n1018 PAR_2_0_VDD075CPU 5.86156794248e-10
L_6_176 PAR_0_3_VDD075CPU n1019 9.3589323149e-08
R_6_176 n1019 PAR_2_0_VDD075CPU 9.87286382756
R_7_176 PAR_0_3_VDD075CPU n1020 162.509895295
C_7_176 n1020 PAR_2_0_VDD075CPU 1.26164578267e-09
G0_177 PAR_0_3_VDD075CPU PAR_0_1_VSS PAR_0_3_VDD075CPU PAR_0_1_VSS -0.748129310261
C0_177 PAR_0_3_VDD075CPU PAR_0_1_VSS 1.65193232601e-10
R_1_177 PAR_0_3_VDD075CPU n1021 0.113290960851
C_1_177 n1021 PAR_0_1_VSS 2.48836096933e-10
R_2_177 PAR_0_3_VDD075CPU n1022 0.461246201526
C_2_177 n1022 PAR_0_1_VSS 2.14228046345e-10
L_3_177 PAR_0_3_VDD075CPU n1023 4.91048903019e-10
R_3_177 n1023 PAR_0_1_VSS 1.52088049943
L_4_177 PAR_0_3_VDD075CPU n1024 7.9487875969e-09
R_4_177 n1024 PAR_0_1_VSS 11.0356447037
R_5_177 PAR_0_3_VDD075CPU n1025 31.2198937002
C_5_177 n1025 PAR_0_1_VSS 2.56697956709e-10
G0_178 PAR_0_3_VDD075CPU PAR_0_1_VDD075CPU PAR_0_3_VDD075CPU PAR_0_1_VDD075CPU -8.35300475006
C0_178 PAR_0_3_VDD075CPU PAR_0_1_VDD075CPU 9.91524620606e-11
R_1_178 PAR_0_3_VDD075CPU n1026 0.4347938192
C_1_178 n1026 PAR_0_1_VDD075CPU 1.10083306467e-10
L_2_178 PAR_0_3_VDD075CPU n1027 2.29152776539e-11
R_2_178 n1027 PAR_0_1_VDD075CPU 0.174401585907
R_3_178 PAR_0_3_VDD075CPU n1028 0.18937688122
C_3_178 n1028 PAR_0_1_VDD075CPU 1.12575909116e-09
L_4_178 PAR_0_3_VDD075CPU n1029 1.75075160611e-10
R_4_178 n1029 PAR_0_1_VDD075CPU 0.426104108181
R_5_178 PAR_0_3_VDD075CPU n1030 1.37952341278
C_5_178 n1030 PAR_0_1_VDD075CPU 8.18342405282e-10
L_6_178 PAR_0_3_VDD075CPU n1031 1.31752793747e-08
R_6_178 n1031 PAR_0_1_VDD075CPU 3.67120728558
R_7_178 PAR_0_3_VDD075CPU n1032 20.9641710715
C_7_178 n1032 PAR_0_1_VDD075CPU 6.48419636692e-10
G0_179 PAR_0_3_VDD075CPU PAR_1_1_VSS PAR_0_3_VDD075CPU PAR_1_1_VSS -3.17196722623
C0_179 PAR_0_3_VDD075CPU PAR_1_1_VSS 8.31678786085e-11
R_1_179 PAR_0_3_VDD075CPU n1033 0.40996391878
C_1_179 n1033 PAR_1_1_VSS 4.72035233235e-11
L_2_179 PAR_0_3_VDD075CPU n1034 1.84513997488e-11
R_2_179 n1034 PAR_1_1_VSS 0.384226890658
R_3_179 PAR_0_3_VDD075CPU n1035 1.96907777459
C_3_179 n1035 PAR_1_1_VSS 6.46911101775e-11
L_4_179 PAR_0_3_VDD075CPU n1036 4.82995312591e-10
R_4_179 n1036 PAR_1_1_VSS 2.03657997297
R_5_179 PAR_0_3_VDD075CPU n1037 4.94417396806
C_5_179 n1037 PAR_1_1_VSS 9.58596619235e-11
L_6_179 PAR_0_3_VDD075CPU n1038 1.76749280147e-08
R_6_179 n1038 PAR_1_1_VSS 13.9585254783
R_7_179 PAR_0_3_VDD075CPU n1039 44.2126440434
C_7_179 n1039 PAR_1_1_VSS 8.85300849998e-11
L_8_179 PAR_0_3_VDD075CPU n1040 2.10304874308e-06
R_8_179 n1040 PAR_1_1_VSS 149.739044225
G0_180 PAR_0_3_VDD075CPU PAR_1_1_VDD075CPU PAR_0_3_VDD075CPU PAR_1_1_VDD075CPU -2.64572486153
C0_180 PAR_0_3_VDD075CPU PAR_1_1_VDD075CPU 9.06841224361e-11
R_1_180 PAR_0_3_VDD075CPU n1041 0.425198029236
C_1_180 n1041 PAR_1_1_VDD075CPU 5.25338205089e-11
L_2_180 PAR_0_3_VDD075CPU n1042 2.15498304158e-11
R_2_180 n1042 PAR_1_1_VDD075CPU 0.421465895007
R_3_180 PAR_0_3_VDD075CPU n1043 4.83989317441
C_3_180 n1043 PAR_1_1_VDD075CPU 2.8536539749e-11
L_4_180 PAR_0_3_VDD075CPU n1044 1.26979675663e-09
R_4_180 n1044 PAR_1_1_VDD075CPU 4.16015493523
R_5_180 PAR_0_3_VDD075CPU n1045 12.1367347586
C_5_180 n1045 PAR_1_1_VDD075CPU 6.59477896411e-11
L_6_180 PAR_0_3_VDD075CPU n1046 8.6439330904e-08
R_6_180 n1046 PAR_1_1_VDD075CPU 30.8578890963
R_7_180 PAR_0_3_VDD075CPU n1047 205.384552122
C_7_180 n1047 PAR_1_1_VDD075CPU 6.1108070969e-11
G0_181 PAR_0_3_VDD075CPU PAR_2_1_VSS PAR_0_3_VDD075CPU PAR_2_1_VSS -2.99092156366
C0_181 PAR_0_3_VDD075CPU PAR_2_1_VSS 1.28367330664e-10
R_1_181 PAR_0_3_VDD075CPU n1048 1.31183952182
C_1_181 n1048 PAR_2_1_VSS 3.86424293699e-11
L_2_181 PAR_0_3_VDD075CPU n1049 6.49906935256e-11
R_2_181 n1049 PAR_2_1_VSS 0.487232973637
R_3_181 PAR_0_3_VDD075CPU n1050 0.51939230768
C_3_181 n1050 PAR_2_1_VSS 3.91843585134e-10
L_4_181 PAR_0_3_VDD075CPU n1051 5.68034874531e-10
R_4_181 n1051 PAR_2_1_VSS 1.2225158552
R_5_181 PAR_0_3_VDD075CPU n1052 3.54168817784
C_5_181 n1052 PAR_2_1_VSS 3.51830852539e-10
L_6_181 PAR_0_3_VDD075CPU n1053 3.34064174256e-08
R_6_181 n1053 PAR_2_1_VSS 8.2966885415
R_7_181 PAR_0_3_VDD075CPU n1054 47.7212158582
C_7_181 n1054 PAR_2_1_VSS 2.9440208042e-10
G0_182 PAR_0_3_VDD075CPU PAR_2_1_VDD075CPU PAR_0_3_VDD075CPU PAR_2_1_VDD075CPU -2.4912755235
C0_182 PAR_0_3_VDD075CPU PAR_2_1_VDD075CPU 9.09716253926e-11
R_1_182 PAR_0_3_VDD075CPU n1055 0.70386227904
C_1_182 n1055 PAR_2_1_VDD075CPU 6.29422345895e-11
L_2_182 PAR_0_3_VDD075CPU n1056 7.01772368119e-11
R_2_182 n1056 PAR_2_1_VDD075CPU 0.512357438502
R_3_182 PAR_0_3_VDD075CPU n1057 1.14708264613
C_3_182 n1057 PAR_2_1_VDD075CPU 3.13154042783e-10
L_4_182 PAR_0_3_VDD075CPU n1058 2.46151539432e-09
R_4_182 n1058 PAR_2_1_VDD075CPU 2.14642339795
R_5_182 PAR_0_3_VDD075CPU n1059 5.03103446547
C_5_182 n1059 PAR_2_1_VDD075CPU 8.95118918647e-10
L_6_182 PAR_0_3_VDD075CPU n1060 2.09000913769e-07
R_6_182 n1060 PAR_2_1_VDD075CPU 13.5842895228
C0_183 PAR_0_3_VDD075CPU PAR_0_2_VSS 1.45490701062e-10
R_1_183 PAR_0_3_VDD075CPU n1061 0.0262580465612
C_1_183 n1061 PAR_0_2_VSS 1.2998104593e-09
R_2_183 PAR_0_3_VDD075CPU n1062 0.151199994141
C_2_183 n1062 PAR_0_2_VSS 3.71368138355e-10
R_3_183 PAR_0_3_VDD075CPU n1063 1.69743365424
C_3_183 n1063 PAR_0_2_VSS 1.02528479188e-10
R_4_183 PAR_0_3_VDD075CPU n1064 17.7539417209
C_4_183 n1064 PAR_0_2_VSS 3.99701167432e-11
R_5_183 PAR_0_3_VDD075CPU n1065 27.2259108919
C_5_183 n1065 PAR_0_2_VSS 1.19574388362e-10
R_6_183 PAR_0_3_VDD075CPU n1066 51.4778987346
C_6_183 n1066 PAR_0_2_VSS 2.31841410639e-10
R0_184 PAR_0_3_VDD075CPU PAR_0_2_VDD075CPU 0.00821422136485
C0_184 PAR_0_3_VDD075CPU PAR_0_2_VDD075CPU 8.34772665482e-11
L_1_184 PAR_0_3_VDD075CPU n1067 7.39282791662e-13
R_1_184 n1067 PAR_0_2_VDD075CPU 0.0348947713135
L_2_184 PAR_0_3_VDD075CPU n1068 7.93401301502e-13
R_2_184 n1068 PAR_0_2_VDD075CPU 0.0203365568695
L_3_184 PAR_0_3_VDD075CPU n1069 7.81231076746e-11
R_3_184 n1069 PAR_0_2_VDD075CPU 0.594375613458
L_4_184 PAR_0_3_VDD075CPU n1070 3.81692356023e-09
R_4_184 n1070 PAR_0_2_VDD075CPU 14.0325280921
L_5_184 PAR_0_3_VDD075CPU n1071 2.28859560421e-07
R_5_184 n1071 PAR_0_2_VDD075CPU 217.929288416
L_6_184 PAR_0_3_VDD075CPU n1072 8.70094684338e-06
R_6_184 n1072 PAR_0_2_VDD075CPU 1183.4463351
G0_185 PAR_0_3_VDD075CPU PAR_1_2_VSS PAR_0_3_VDD075CPU PAR_1_2_VSS -0.3345672681
C0_185 PAR_0_3_VDD075CPU PAR_1_2_VSS 1.42023224721e-10
R_1_185 PAR_0_3_VDD075CPU n1073 0.233842948493
C_1_185 n1073 PAR_1_2_VSS 1.37092702446e-10
R_2_185 PAR_0_3_VDD075CPU n1074 3.54930525884
C_2_185 n1074 PAR_1_2_VSS 3.38819444918e-11
L_3_185 PAR_0_3_VDD075CPU n1075 7.84205952823e-10
R_3_185 n1075 PAR_1_2_VSS 3.23959643916
L_4_185 PAR_0_3_VDD075CPU n1076 1.5825902516e-07
R_4_185 n1076 PAR_1_2_VSS 64.9066866849
L_5_185 PAR_0_3_VDD075CPU n1077 9.60118235511e-07
R_5_185 n1077 PAR_1_2_VSS 95.4188095805
R0_186 PAR_0_3_VDD075CPU PAR_1_2_VDD075CPU 0.401482240089
C0_186 PAR_0_3_VDD075CPU PAR_1_2_VDD075CPU 1.57028347009e-10
L_1_186 PAR_0_3_VDD075CPU n1078 8.08542567319e-12
R_1_186 n1078 PAR_1_2_VDD075CPU 0.215832365293
L_2_186 PAR_0_3_VDD075CPU n1079 1.54794746865e-10
R_2_186 n1079 PAR_1_2_VDD075CPU 1.97198902666
L_3_186 PAR_0_3_VDD075CPU n1080 6.60750838077e-10
R_3_186 n1080 PAR_1_2_VDD075CPU 3.9945744578
L_4_186 PAR_0_3_VDD075CPU n1081 4.34787104027e-08
R_4_186 n1081 PAR_1_2_VDD075CPU 77.327314856
L_5_186 PAR_0_3_VDD075CPU n1082 2.87884586301e-06
R_5_186 n1082 PAR_1_2_VDD075CPU 690.057679303
L_6_186 PAR_0_3_VDD075CPU n1083 0.0019656837274
R_6_186 n1083 PAR_1_2_VDD075CPU 4984.50462902
G0_187 PAR_0_3_VDD075CPU PAR_2_2_VSS PAR_0_3_VDD075CPU PAR_2_2_VSS -0.185207159753
C0_187 PAR_0_3_VDD075CPU PAR_2_2_VSS 3.02454387134e-11
R_1_187 PAR_0_3_VDD075CPU n1084 0.17692372962
C_1_187 n1084 PAR_2_2_VSS 1.30838046602e-10
R_2_187 PAR_0_3_VDD075CPU n1085 2.67644402436
C_2_187 n1085 PAR_2_2_VSS 4.35435139987e-11
L_3_187 PAR_0_3_VDD075CPU n1086 2.31007927814e-09
R_3_187 n1086 PAR_2_2_VSS 7.58901880127
L_4_187 PAR_0_3_VDD075CPU n1087 2.24557515017e-08
R_4_187 n1087 PAR_2_2_VSS 27.6732186803
L_5_187 PAR_0_3_VDD075CPU n1088 2.64733699847e-07
R_5_187 n1088 PAR_2_2_VSS 79.7687124828
L_6_187 PAR_0_3_VDD075CPU n1089 2.63494480875e-06
R_6_187 n1089 PAR_2_2_VSS 209.839017454
G0_188 PAR_0_3_VDD075CPU PAR_2_2_VDD075CPU PAR_0_3_VDD075CPU PAR_2_2_VDD075CPU -0.242473928223
C0_188 PAR_0_3_VDD075CPU PAR_2_2_VDD075CPU 1.81214225897e-11
R_1_188 PAR_0_3_VDD075CPU n1090 2.47738324619
C_1_188 n1090 PAR_2_2_VDD075CPU 7.30940599529e-12
L_2_188 PAR_0_3_VDD075CPU n1091 5.07377508395e-10
R_2_188 n1091 PAR_2_2_VDD075CPU 6.84462972648
L_3_188 PAR_0_3_VDD075CPU n1092 1.41225959477e-09
R_3_188 n1092 PAR_2_2_VDD075CPU 10.4737859375
L_4_188 PAR_0_3_VDD075CPU n1093 8.14475860934e-07
R_4_188 n1093 PAR_2_2_VDD075CPU 1319.79193624
L_5_188 PAR_0_3_VDD075CPU n1094 3.71517654885e-05
R_5_188 n1094 PAR_2_2_VDD075CPU 8227.81765351
R_1_189 PAR_0_3_VDD075CPU n1095 0.00067517335272
C_1_189 n1095 PAR_0_3_VSS 2.89028179015e-08
R_2_189 PAR_0_3_VDD075CPU n1096 0.000646920309506
C_2_189 n1096 PAR_0_3_VSS 5.93043808698e-08
R_3_189 PAR_0_3_VDD075CPU n1097 0.0550662979999
C_3_189 n1097 PAR_0_3_VSS 2.58971889822e-09
R_4_189 PAR_0_3_VDD075CPU n1098 0.249642204989
C_4_189 n1098 PAR_0_3_VSS 1.21144285564e-09
R_5_189 PAR_0_3_VDD075CPU n1099 3.84683789549
C_5_189 n1099 PAR_0_3_VSS 2.77907998244e-10
R_6_189 PAR_0_3_VDD075CPU n1100 16.3084281032
C_6_189 n1100 PAR_0_3_VSS 4.36095876241e-10
G0_190 PAR_0_3_VDD075CPU PAR_0_0_VSS PAR_0_3_VDD075CPU PAR_0_0_VSS -2.15709267362
C0_190 PAR_0_3_VDD075CPU PAR_0_0_VSS 2.10783687757e-10
R_1_190 PAR_0_3_VDD075CPU n1101 0.0178014117789
C_1_190 n1101 PAR_0_0_VSS 1.05700404469e-09
R_2_190 PAR_0_3_VDD075CPU n1102 0.844042493521
C_2_190 n1102 PAR_0_0_VSS 1.72486472486e-10
L_3_190 PAR_0_3_VDD075CPU n1103 1.20498378944e-10
R_3_190 n1103 PAR_0_0_VSS 0.482965646938
L_4_190 PAR_0_3_VDD075CPU n1104 8.29293187449e-09
R_4_190 n1104 PAR_0_0_VSS 11.5537432641
R_5_190 PAR_0_3_VDD075CPU n1105 565.926390034
C_5_190 n1105 PAR_0_0_VSS 3.45361092361e-11
G0_191 PAR_1_3_VSS PAR_0_0_VDD075CPU PAR_1_3_VSS PAR_0_0_VDD075CPU -0.0802824274004
C0_191 PAR_1_3_VSS PAR_0_0_VDD075CPU 1.8920135235e-10
R_1_191 PAR_1_3_VSS n1106 0.146329861153
C_1_191 n1106 PAR_0_0_VDD075CPU 2.2993971438e-10
R_2_191 PAR_1_3_VSS n1107 0.430361263849
C_2_191 n1107 PAR_0_0_VDD075CPU 2.20990859953e-10
R_3_191 PAR_1_3_VSS n1108 4.57739679448
C_3_191 n1108 PAR_0_0_VDD075CPU 6.50125672612e-11
R_4_191 PAR_1_3_VSS n1109 10.811107402
C_4_191 n1109 PAR_0_0_VDD075CPU 2.18153334794e-10
L_5_191 PAR_1_3_VSS n1110 9.76858540139e-08
R_5_191 n1110 PAR_0_0_VDD075CPU 12.4560255475
G0_192 PAR_1_3_VSS PAR_1_0_VSS PAR_1_3_VSS PAR_1_0_VSS -0.735103856456
C0_192 PAR_1_3_VSS PAR_1_0_VSS 1.60537338302e-10
R_1_192 PAR_1_3_VSS n1111 0.385136917311
C_1_192 n1111 PAR_1_0_VSS 2.45926434605e-10
R_2_192 PAR_1_3_VSS n1112 0.0867840329915
C_2_192 n1112 PAR_1_0_VSS 3.61340286003e-09
R_3_192 PAR_1_3_VSS n1113 0.150120033109
C_3_192 n1113 PAR_1_0_VSS 8.38209337955e-09
L_4_192 PAR_1_3_VSS n1114 1.68209541221e-08
R_4_192 n1114 PAR_1_0_VSS 1.36029067135
G0_193 PAR_1_3_VSS PAR_1_0_VDD075CPU PAR_1_3_VSS PAR_1_0_VDD075CPU -0.0878379170289
C0_193 PAR_1_3_VSS PAR_1_0_VDD075CPU 1.99787573388e-10
R_1_193 PAR_1_3_VSS n1115 0.178581119819
C_1_193 n1115 PAR_1_0_VDD075CPU 2.16711608786e-10
R_2_193 PAR_1_3_VSS n1116 0.427813870116
C_2_193 n1116 PAR_1_0_VDD075CPU 2.29904831119e-10
R_3_193 PAR_1_3_VSS n1117 3.31129347449
C_3_193 n1117 PAR_1_0_VDD075CPU 8.06983408826e-11
R_4_193 PAR_1_3_VSS n1118 8.38089034972
C_4_193 n1118 PAR_1_0_VDD075CPU 2.76015738438e-10
L_5_193 PAR_1_3_VSS n1119 8.71846884243e-08
R_5_193 n1119 PAR_1_0_VDD075CPU 11.3846047637
G0_194 PAR_1_3_VSS PAR_2_0_VSS PAR_1_3_VSS PAR_2_0_VSS -1.53309104696
C0_194 PAR_1_3_VSS PAR_2_0_VSS 2.11134441076e-10
R_1_194 PAR_1_3_VSS n1120 0.266454294352
C_1_194 n1120 PAR_2_0_VSS 1.87336674931e-10
R_2_194 PAR_1_3_VSS n1121 1.19990975644
C_2_194 n1121 PAR_2_0_VSS 9.05550772579e-11
R_3_194 PAR_1_3_VSS n1122 0.189539890417
C_3_194 n1122 PAR_2_0_VSS 3.73624612237e-09
R_4_194 PAR_1_3_VSS n1123 0.137322840383
C_4_194 n1123 PAR_2_0_VSS 1.13810787358e-08
L_5_194 PAR_1_3_VSS n1124 4.42354153627e-09
R_5_194 n1124 PAR_2_0_VSS 0.89710728706
L_6_194 PAR_1_3_VSS n1125 3.54028282521e-08
R_6_194 n1125 PAR_2_0_VSS 2.39007015465
G0_195 PAR_1_3_VSS PAR_2_0_VDD075CPU PAR_1_3_VSS PAR_2_0_VDD075CPU -0.0946822409661
C0_195 PAR_1_3_VSS PAR_2_0_VDD075CPU 2.09331801671e-10
R_1_195 PAR_1_3_VSS n1126 0.168704463135
C_1_195 n1126 PAR_2_0_VDD075CPU 2.12651422256e-10
R_2_195 PAR_1_3_VSS n1127 0.369349567743
C_2_195 n1127 PAR_2_0_VDD075CPU 2.49710261537e-10
R_3_195 PAR_1_3_VSS n1128 1.31296060812
C_3_195 n1128 PAR_2_0_VDD075CPU 1.91851833603e-10
R_4_195 PAR_1_3_VSS n1129 7.82196170721
C_4_195 n1129 PAR_2_0_VDD075CPU 2.77271450043e-10
L_5_195 PAR_1_3_VSS n1130 8.46825515344e-08
R_5_195 n1130 PAR_2_0_VDD075CPU 10.561642403
R0_196 PAR_1_3_VSS PAR_0_1_VSS 99.5332185535
C0_196 PAR_1_3_VSS PAR_0_1_VSS 1.14089881752e-10
R_1_196 PAR_1_3_VSS n1131 0.23238450857
C_1_196 n1131 PAR_0_1_VSS 5.12154208641e-10
R_2_196 PAR_1_3_VSS n1132 0.0886453632787
C_2_196 n1132 PAR_0_1_VSS 3.76575240092e-09
R_3_196 PAR_1_3_VSS n1133 0.289122655757
C_3_196 n1133 PAR_0_1_VSS 2.94545675799e-09
R_4_196 PAR_1_3_VSS n1134 0.19054085571
C_4_196 n1134 PAR_0_1_VSS 1.76986468044e-08
R_5_196 PAR_1_3_VSS n1135 0.714533049455
C_5_196 n1135 PAR_0_1_VSS 1.82725388262e-08
G0_197 PAR_1_3_VSS PAR_0_1_VDD075CPU PAR_1_3_VSS PAR_0_1_VDD075CPU -0.0676683020442
C0_197 PAR_1_3_VSS PAR_0_1_VDD075CPU 1.53450572312e-10
R_1_197 PAR_1_3_VSS n1136 0.198552173517
C_1_197 n1136 PAR_0_1_VDD075CPU 1.81047115329e-10
R_2_197 PAR_1_3_VSS n1137 0.629386127638
C_2_197 n1137 PAR_0_1_VDD075CPU 1.46993234079e-10
R_3_197 PAR_1_3_VSS n1138 2.52079642254
C_3_197 n1138 PAR_0_1_VDD075CPU 9.864600114e-11
R_4_197 PAR_1_3_VSS n1139 9.18311499236
C_4_197 n1139 PAR_0_1_VDD075CPU 2.18444630578e-10
L_5_197 PAR_1_3_VSS n1140 1.16337182917e-07
R_5_197 n1140 PAR_0_1_VDD075CPU 14.7779673718
G0_198 PAR_1_3_VSS PAR_1_1_VSS PAR_1_3_VSS PAR_1_1_VSS -0.0367220833258
C0_198 PAR_1_3_VSS PAR_1_1_VSS 1.24225972154e-10
R_1_198 PAR_1_3_VSS n1141 0.31454937561
C_1_198 n1141 PAR_1_1_VSS 1.1573458894e-10
R_2_198 PAR_1_3_VSS n1142 3.89436820043
C_2_198 n1142 PAR_1_1_VSS 2.87538540821e-11
R_3_198 PAR_1_3_VSS n1143 4.54448694863
C_3_198 n1143 PAR_1_1_VSS 6.40262654352e-11
R_4_198 PAR_1_3_VSS n1144 14.8163572025
C_4_198 n1144 PAR_1_1_VSS 1.3029340783e-10
L_5_198 PAR_1_3_VSS n1145 2.06400996062e-07
R_5_198 n1145 PAR_1_1_VSS 25.8370162202
G0_199 PAR_1_3_VSS PAR_1_1_VDD075CPU PAR_1_3_VSS PAR_1_1_VDD075CPU -0.0458489744278
C0_199 PAR_1_3_VSS PAR_1_1_VDD075CPU 1.29526986899e-10
R_1_199 PAR_1_3_VSS n1146 0.291731195745
C_1_199 n1146 PAR_1_1_VDD075CPU 1.21329153207e-10
R_2_199 PAR_1_3_VSS n1147 1.22990749965
C_2_199 n1147 PAR_1_1_VDD075CPU 7.25458181551e-11
R_3_199 PAR_1_3_VSS n1148 2.81561021617
C_3_199 n1148 PAR_1_1_VDD075CPU 9.30946711852e-11
R_4_199 PAR_1_3_VSS n1149 11.3124665628
C_4_199 n1149 PAR_1_1_VDD075CPU 1.5998101083e-10
L_5_199 PAR_1_3_VSS n1150 1.8095676939e-07
R_5_199 n1150 PAR_1_1_VDD075CPU 21.8107374234
R0_200 PAR_1_3_VSS PAR_2_1_VSS 2.49963126697
C0_200 PAR_1_3_VSS PAR_2_1_VSS 1.57081504827e-10
R_1_200 PAR_1_3_VSS n1151 0.276906799635
C_1_200 n1151 PAR_2_1_VSS 1.33958954092e-10
R_2_200 PAR_1_3_VSS n1152 1.8129342286
C_2_200 n1152 PAR_2_1_VSS 1.06883711383e-10
R_3_200 PAR_1_3_VSS n1153 0.271675594089
C_3_200 n1153 PAR_2_1_VSS 1.59317307664e-09
L_4_200 PAR_1_3_VSS n1154 4.04455846438e-09
R_4_200 n1154 PAR_2_1_VSS 2.60712263713
L_5_200 PAR_1_3_VSS n1155 8.08127425436e-09
R_5_200 n1155 PAR_2_1_VSS 1.8814671179
L_6_200 PAR_1_3_VSS n1156 1.022646296e-07
R_6_200 n1156 PAR_2_1_VSS 7.07350099665
G0_201 PAR_1_3_VSS PAR_2_1_VDD075CPU PAR_1_3_VSS PAR_2_1_VDD075CPU -0.0557780995941
C0_201 PAR_1_3_VSS PAR_2_1_VDD075CPU 1.52349526234e-10
R_1_201 PAR_1_3_VSS n1157 0.230729114111
C_1_201 n1157 PAR_2_1_VDD075CPU 1.96591694533e-10
R_2_201 PAR_1_3_VSS n1158 0.63899072508
C_2_201 n1158 PAR_2_1_VDD075CPU 2.0505013255e-10
R_3_201 PAR_1_3_VSS n1159 11.3637114864
C_3_201 n1159 PAR_2_1_VDD075CPU 2.8149551039e-10
L_4_201 PAR_1_3_VSS n1160 2.52303492861e-07
R_4_201 n1160 PAR_2_1_VDD075CPU 17.9281825426
R0_202 PAR_1_3_VSS PAR_0_2_VSS 0.508940399129
C0_202 PAR_1_3_VSS PAR_0_2_VSS 1.48995898452e-10
L_1_202 PAR_1_3_VSS n1161 4.24239818794e-12
R_1_202 n1161 PAR_0_2_VSS 0.165047859328
R_2_202 PAR_1_3_VSS n1162 0.173084762147
C_2_202 n1162 PAR_0_2_VSS 7.60615731882e-10
R_3_202 PAR_1_3_VSS n1163 0.0992516018258
C_3_202 n1163 PAR_0_2_VSS 3.96866096203e-09
R_4_202 PAR_1_3_VSS n1164 0.398846754279
C_4_202 n1164 PAR_0_2_VSS 3.30696470664e-09
R_5_202 PAR_1_3_VSS n1165 0.22474385364
C_5_202 n1165 PAR_0_2_VSS 1.70229520096e-08
R_6_202 PAR_1_3_VSS n1166 0.849802720883
C_6_202 n1166 PAR_0_2_VSS 1.58027450735e-08
G0_203 PAR_1_3_VSS PAR_0_2_VDD075CPU PAR_1_3_VSS PAR_0_2_VDD075CPU -0.232604466056
C0_203 PAR_1_3_VSS PAR_0_2_VDD075CPU 1.75891010843e-10
R_1_203 PAR_1_3_VSS n1167 0.100399709687
C_1_203 n1167 PAR_0_2_VDD075CPU 3.92869794442e-10
R_2_203 PAR_1_3_VSS n1168 0.809896028577
C_2_203 n1168 PAR_0_2_VDD075CPU 1.50864767761e-10
R_3_203 PAR_1_3_VSS n1169 12.0602709157
C_3_203 n1169 PAR_0_2_VDD075CPU 3.78479150635e-11
R_4_203 PAR_1_3_VSS n1170 4.12402787717
C_4_203 n1170 PAR_0_2_VDD075CPU 9.20598250896e-10
L_5_203 PAR_1_3_VSS n1171 2.32950683197e-08
R_5_203 n1171 PAR_0_2_VDD075CPU 4.29914354089
R0_204 PAR_1_3_VSS PAR_1_2_VSS 0.00746474964779
C0_204 PAR_1_3_VSS PAR_1_2_VSS 6.15999751368e-11
L_1_204 PAR_1_3_VSS n1172 5.6203216904e-13
R_1_204 n1172 PAR_1_2_VSS 0.0138839187466
L_2_204 PAR_1_3_VSS n1173 5.61601389798e-11
R_2_204 n1173 PAR_1_2_VSS 0.245147825508
R_3_204 PAR_1_3_VSS n1174 0.537114122663
C_3_204 n1174 PAR_1_2_VSS 1.00977628809e-09
L_4_204 PAR_1_3_VSS n1175 3.01946214941e-10
R_4_204 n1175 PAR_1_2_VSS 0.157136123213
L_5_204 PAR_1_3_VSS n1176 6.31916838156e-09
R_5_204 n1176 PAR_1_2_VSS 0.778196400278
G0_205 PAR_1_3_VSS PAR_1_2_VDD075CPU PAR_1_3_VSS PAR_1_2_VDD075CPU -0.0607220865784
C0_205 PAR_1_3_VSS PAR_1_2_VDD075CPU 1.80126944448e-10
R_1_205 PAR_1_3_VSS n1177 0.0100391478389
C_1_205 n1177 PAR_1_2_VDD075CPU 2.95941914493e-09
R_2_205 PAR_1_3_VSS n1178 0.0198635099975
C_2_205 n1178 PAR_1_2_VDD075CPU 2.31793371918e-09
R_3_205 PAR_1_3_VSS n1179 1.36343450947
C_3_205 n1179 PAR_1_2_VDD075CPU 1.68718004536e-10
R_4_205 PAR_1_3_VSS n1180 7.33231099596
C_4_205 n1180 PAR_1_2_VDD075CPU 2.38280499667e-10
L_5_205 PAR_1_3_VSS n1181 1.416935327e-07
R_5_205 n1181 PAR_1_2_VDD075CPU 16.4684716639
R0_206 PAR_1_3_VSS PAR_2_2_VSS 0.638390545383
C0_206 PAR_1_3_VSS PAR_2_2_VSS 1.70072110719e-11
R_1_206 PAR_1_3_VSS n1182 0.307736282051
C_1_206 n1182 PAR_2_2_VSS 2.86156522617e-10
R_2_206 PAR_1_3_VSS n1183 0.200959783867
C_2_206 n1183 PAR_2_2_VSS 2.43250477132e-09
L_3_206 PAR_1_3_VSS n1184 7.09879739995e-10
R_3_206 n1184 PAR_2_2_VSS 0.452098011273
L_4_206 PAR_1_3_VSS n1185 3.1983527778e-09
R_4_206 n1185 PAR_2_2_VSS 0.771947257762
L_5_206 PAR_1_3_VSS n1186 4.91206884598e-08
R_5_206 n1186 PAR_2_2_VSS 3.41535864614
C0_207 PAR_1_3_VSS PAR_2_2_VDD075CPU 2.09415525882e-11
R_1_207 PAR_1_3_VSS n1187 0.835288460953
C_1_207 n1187 PAR_2_2_VDD075CPU 7.38732231836e-11
R_2_207 PAR_1_3_VSS n1188 1315.03560416
C_2_207 n1188 PAR_2_2_VDD075CPU 1.60790924498e-11
R0_208 PAR_1_3_VSS PAR_0_3_VSS 0.00439652877915
L_1_208 PAR_1_3_VSS n1189 3.09384003233e-13
R_1_208 n1189 PAR_0_3_VSS 0.00977685518214
R_2_208 PAR_1_3_VSS n1190 0.0645466623715
C_2_208 n1190 PAR_0_3_VSS 4.52450366289e-09
L_3_208 PAR_1_3_VSS n1191 7.22682656568e-11
R_3_208 n1191 PAR_0_3_VSS 0.143571866495
R_4_208 PAR_1_3_VSS n1192 0.139720331085
C_4_208 n1192 PAR_0_3_VSS 1.44988852421e-08
R_5_208 PAR_1_3_VSS n1193 0.293428262387
C_5_208 n1193 PAR_0_3_VSS 1.6561955315e-08
R_6_208 PAR_1_3_VSS n1194 1.0000230122
C_6_208 n1194 PAR_0_3_VSS 1.46285103779e-08
G0_209 PAR_1_3_VSS PAR_0_3_VDD075CPU PAR_1_3_VSS PAR_0_3_VDD075CPU -0.0318487916914
C0_209 PAR_1_3_VSS PAR_0_3_VDD075CPU 1.39375999235e-10
R_1_209 PAR_1_3_VSS n1195 0.0148250614851
C_1_209 n1195 PAR_0_3_VDD075CPU 2.24760422187e-09
R_2_209 PAR_1_3_VSS n1196 0.265147127284
C_2_209 n1196 PAR_0_3_VDD075CPU 3.46323509887e-10
L_3_209 PAR_1_3_VSS n1197 4.00951022414e-07
R_3_209 n1197 PAR_0_3_VDD075CPU 331.133411008
L_4_209 PAR_1_3_VSS n1198 3.22784647853e-07
R_4_209 n1198 PAR_0_3_VDD075CPU 34.6874581126
R0_210 PAR_1_3_VSS PAR_0_0_VSS 126.454410783
C0_210 PAR_1_3_VSS PAR_0_0_VSS 1.63724356156e-10
R_1_210 PAR_1_3_VSS n1199 0.0357771923235
C_1_210 n1199 PAR_0_0_VSS 1.54073206094e-09
R_2_210 PAR_1_3_VSS n1200 0.0775200070694
C_2_210 n1200 PAR_0_0_VSS 1.83485270436e-09
R_3_210 PAR_1_3_VSS n1201 0.0568857053181
C_3_210 n1201 PAR_0_0_VSS 6.41825534797e-09
R_4_210 PAR_1_3_VSS n1202 0.188315006209
C_4_210 n1202 PAR_0_0_VSS 6.68116243478e-09
R_5_210 PAR_1_3_VSS n1203 0.0626935740551
C_5_210 n1203 PAR_0_0_VSS 4.01445201806e-08
R_6_210 PAR_1_3_VSS n1204 1.84276337478
C_6_210 n1204 PAR_0_0_VSS 6.78994965234e-09
G0_211 PAR_1_3_VDD075CPU PAR_0_0_VDD075CPU PAR_1_3_VDD075CPU PAR_0_0_VDD075CPU -6.76022723786
C0_211 PAR_1_3_VDD075CPU PAR_0_0_VDD075CPU 1.167749708e-10
R_1_211 PAR_1_3_VDD075CPU n1205 0.280959572497
C_1_211 n1205 PAR_0_0_VDD075CPU 1.34004837716e-10
L_2_211 PAR_1_3_VDD075CPU n1206 1.50501699091e-11
R_2_211 n1206 PAR_0_0_VDD075CPU 0.178819283693
R_3_211 PAR_1_3_VDD075CPU n1207 0.359484847758
C_3_211 n1207 PAR_0_0_VDD075CPU 4.1864071567e-10
L_4_211 PAR_1_3_VDD075CPU n1208 3.60518675956e-10
R_4_211 n1208 PAR_0_0_VDD075CPU 1.00996657524
R_5_211 PAR_1_3_VDD075CPU n1209 2.53170955554
C_5_211 n1209 PAR_0_0_VDD075CPU 4.13151598252e-10
L_6_211 PAR_1_3_VDD075CPU n1210 1.67145415977e-08
R_6_211 n1210 PAR_0_0_VDD075CPU 5.6185255675
R_7_211 PAR_1_3_VDD075CPU n1211 41.2407209752
C_7_211 n1211 PAR_0_0_VDD075CPU 3.23353189027e-10
G0_212 PAR_1_3_VDD075CPU PAR_1_0_VSS PAR_1_3_VDD075CPU PAR_1_0_VSS -0.405138231726
C0_212 PAR_1_3_VDD075CPU PAR_1_0_VSS 1.6335130063e-10
R_1_212 PAR_1_3_VDD075CPU n1212 0.199985304206
C_1_212 n1212 PAR_1_0_VSS 1.43026325017e-10
R_2_212 PAR_1_3_VDD075CPU n1213 1.85073934605
C_2_212 n1213 PAR_1_0_VSS 6.01621834139e-11
L_3_212 PAR_1_3_VDD075CPU n1214 1.02431847558e-09
R_3_212 n1214 PAR_1_0_VSS 3.03404971765
L_4_212 PAR_1_3_VDD075CPU n1215 2.42284142731e-08
R_4_212 n1215 PAR_1_0_VSS 15.1323821405
L_5_212 PAR_1_3_VDD075CPU n1216 9.7384860015e-07
R_5_212 n1216 PAR_1_0_VSS 107.664582456
L_6_212 PAR_1_3_VDD075CPU n1217 0.00130229917278
R_6_212 n1217 PAR_1_0_VSS 5740.84874774
G0_213 PAR_1_3_VDD075CPU PAR_1_0_VDD075CPU PAR_1_3_VDD075CPU PAR_1_0_VDD075CPU -4.42299741746
C0_213 PAR_1_3_VDD075CPU PAR_1_0_VDD075CPU 1.30949751448e-10
R_1_213 PAR_1_3_VDD075CPU n1218 0.326608459244
C_1_213 n1218 PAR_1_0_VDD075CPU 6.96817185086e-11
L_2_213 PAR_1_3_VDD075CPU n1219 1.6565340854e-11
R_2_213 n1219 PAR_1_0_VDD075CPU 0.275404600941
R_3_213 PAR_1_3_VDD075CPU n1220 0.985881789923
C_3_213 n1220 PAR_1_0_VDD075CPU 1.18456989191e-10
L_4_213 PAR_1_3_VDD075CPU n1221 3.94578299317e-10
R_4_213 n1221 PAR_1_0_VDD075CPU 1.49225139452
R_5_213 PAR_1_3_VDD075CPU n1222 3.26327627585
C_5_213 n1222 PAR_1_0_VDD075CPU 1.59645633825e-10
L_6_213 PAR_1_3_VDD075CPU n1223 1.43048930684e-08
R_6_213 n1223 PAR_1_0_VDD075CPU 9.19671429193
R_7_213 PAR_1_3_VDD075CPU n1224 24.7118114834
C_7_213 n1224 PAR_1_0_VDD075CPU 1.960148206e-10
L_8_213 PAR_1_3_VDD075CPU n1225 1.17995104664e-06
R_8_213 n1225 PAR_1_0_VDD075CPU 76.9450682322
G0_214 PAR_1_3_VDD075CPU PAR_2_0_VSS PAR_1_3_VDD075CPU PAR_2_0_VSS -0.431252454154
C0_214 PAR_1_3_VDD075CPU PAR_2_0_VSS 1.89450646432e-10
R_1_214 PAR_1_3_VDD075CPU n1226 0.703199013995
C_1_214 n1226 PAR_2_0_VSS 3.93676711736e-11
L_2_214 PAR_1_3_VDD075CPU n1227 2.49204111163e-10
R_2_214 n1227 PAR_2_0_VSS 2.90188668848
R_3_214 PAR_1_3_VDD075CPU n1228 5.45075274918
C_3_214 n1228 PAR_2_0_VSS 2.82668495503e-11
R_4_214 PAR_1_3_VDD075CPU n1229 7.60730881705
C_4_214 n1229 PAR_2_0_VSS 6.36408276295e-11
L_5_214 PAR_1_3_VDD075CPU n1230 2.27847116638e-08
R_5_214 n1230 PAR_2_0_VSS 12.8338162283
L_6_214 PAR_1_3_VDD075CPU n1231 1.25693151443e-06
R_6_214 n1231 PAR_2_0_VSS 114.548622132
G0_215 PAR_1_3_VDD075CPU PAR_2_0_VDD075CPU PAR_1_3_VDD075CPU PAR_2_0_VDD075CPU -4.18510622162
C0_215 PAR_1_3_VDD075CPU PAR_2_0_VDD075CPU 1.41902127468e-10
R_1_215 PAR_1_3_VDD075CPU n1232 0.309609636223
C_1_215 n1232 PAR_2_0_VDD075CPU 7.541624356e-11
L_2_215 PAR_1_3_VDD075CPU n1233 1.62978514238e-11
R_2_215 n1233 PAR_2_0_VDD075CPU 0.277747807969
R_3_215 PAR_1_3_VDD075CPU n1234 1.36866213452
C_3_215 n1234 PAR_2_0_VDD075CPU 8.79708667361e-11
L_4_215 PAR_1_3_VDD075CPU n1235 5.63872995928e-10
R_4_215 n1235 PAR_2_0_VDD075CPU 1.93916161568
R_5_215 PAR_1_3_VDD075CPU n1236 4.703092467
C_5_215 n1236 PAR_2_0_VDD075CPU 1.2828529054e-10
L_6_215 PAR_1_3_VDD075CPU n1237 2.98337908633e-08
R_6_215 n1237 PAR_2_0_VDD075CPU 15.2960614383
R_7_215 PAR_1_3_VDD075CPU n1238 83.5699414678
C_7_215 n1238 PAR_2_0_VDD075CPU 1.21553918677e-10
L_8_215 PAR_1_3_VDD075CPU n1239 2.29695103036e-05
R_8_215 n1239 PAR_2_0_VDD075CPU 274.328016949
G0_216 PAR_1_3_VDD075CPU PAR_0_1_VSS PAR_1_3_VDD075CPU PAR_0_1_VSS -0.2423650587
C0_216 PAR_1_3_VDD075CPU PAR_0_1_VSS 1.59192563975e-10
R_1_216 PAR_1_3_VDD075CPU n1240 0.139667595161
C_1_216 n1240 PAR_0_1_VSS 1.97805002414e-10
R_2_216 PAR_1_3_VDD075CPU n1241 0.797648775411
C_2_216 n1241 PAR_0_1_VSS 8.04259651492e-11
L_3_216 PAR_1_3_VDD075CPU n1242 1.86224427813e-09
R_3_216 n1242 PAR_0_1_VSS 4.12600724927
R_4_216 PAR_1_3_VDD075CPU n1243 36.9879979105
C_4_216 n1243 PAR_0_1_VSS 2.44364076202e-10
G0_217 PAR_1_3_VDD075CPU PAR_0_1_VDD075CPU PAR_1_3_VDD075CPU PAR_0_1_VDD075CPU -4.19772610484
C0_217 PAR_1_3_VDD075CPU PAR_0_1_VDD075CPU 1.02009393901e-10
R_1_217 PAR_1_3_VDD075CPU n1244 0.309220624397
C_1_217 n1244 PAR_0_1_VDD075CPU 9.19329119435e-11
L_2_217 PAR_1_3_VDD075CPU n1245 1.54678444188e-11
R_2_217 n1245 PAR_0_1_VDD075CPU 0.269285576986
R_3_217 PAR_1_3_VDD075CPU n1246 1.28939674824
C_3_217 n1246 PAR_0_1_VDD075CPU 9.36864278113e-11
L_4_217 PAR_1_3_VDD075CPU n1247 7.01357443433e-10
R_4_217 n1247 PAR_0_1_VDD075CPU 2.35712348311
R_5_217 PAR_1_3_VDD075CPU n1248 5.49066140705
C_5_217 n1248 PAR_0_1_VDD075CPU 1.20382851101e-10
L_6_217 PAR_1_3_VDD075CPU n1249 3.32778427136e-08
R_6_217 n1249 PAR_0_1_VDD075CPU 16.7341080488
R_7_217 PAR_1_3_VDD075CPU n1250 163.793019664
C_7_217 n1250 PAR_0_1_VDD075CPU 6.66151336268e-11
G0_218 PAR_1_3_VDD075CPU PAR_1_1_VSS PAR_1_3_VDD075CPU PAR_1_1_VSS -3.48709236
C0_218 PAR_1_3_VDD075CPU PAR_1_1_VSS 7.91799171317e-11
R_1_218 PAR_1_3_VDD075CPU n1251 0.42087130552
C_1_218 n1251 PAR_1_1_VSS 3.14625354888e-11
L_2_218 PAR_1_3_VDD075CPU n1252 1.48152160614e-11
R_2_218 n1252 PAR_1_1_VSS 0.337366766724
R_3_218 PAR_1_3_VDD075CPU n1253 1.09682654829
C_3_218 n1253 PAR_1_1_VSS 7.03676841092e-11
L_4_218 PAR_1_3_VDD075CPU n1254 3.72119867362e-10
R_4_218 n1254 PAR_1_1_VSS 2.41088313391
R_5_218 PAR_1_3_VDD075CPU n1255 6.09695592033
C_5_218 n1255 PAR_1_1_VSS 5.39681854823e-11
L_6_218 PAR_1_3_VDD075CPU n1256 6.67898832016e-09
R_6_218 n1256 PAR_1_1_VSS 10.4419601771
R_7_218 PAR_1_3_VDD075CPU n1257 29.5885745328
C_7_218 n1257 PAR_1_1_VSS 5.14707607079e-11
L_8_218 PAR_1_3_VDD075CPU n1258 3.24538154758e-07
R_8_218 n1258 PAR_1_1_VSS 80.6058984865
R_9_218 PAR_1_3_VDD075CPU n1259 651.534572236
C_9_218 n1259 PAR_1_1_VSS 2.18765953984e-11
G0_219 PAR_1_3_VDD075CPU PAR_1_1_VDD075CPU PAR_1_3_VDD075CPU PAR_1_1_VDD075CPU -2.6659855136
C0_219 PAR_1_3_VDD075CPU PAR_1_1_VDD075CPU 8.53257297157e-11
R_1_219 PAR_1_3_VDD075CPU n1260 0.491556558623
C_1_219 n1260 PAR_1_1_VDD075CPU 2.89125148234e-11
L_2_219 PAR_1_3_VDD075CPU n1261 2.14414234657e-11
R_2_219 n1261 PAR_1_1_VDD075CPU 0.439544928118
R_3_219 PAR_1_3_VDD075CPU n1262 1.96664939807
C_3_219 n1262 PAR_1_1_VDD075CPU 5.03786162376e-11
L_4_219 PAR_1_3_VDD075CPU n1263 5.69160532012e-10
R_4_219 n1263 PAR_1_1_VDD075CPU 2.88828321342
R_5_219 PAR_1_3_VDD075CPU n1264 9.16978414915
C_5_219 n1264 PAR_1_1_VDD075CPU 4.28581479347e-11
L_6_219 PAR_1_3_VDD075CPU n1265 2.88576220946e-08
R_6_219 n1265 PAR_1_1_VDD075CPU 24.5117861555
R_7_219 PAR_1_3_VDD075CPU n1266 70.9282448385
C_7_219 n1266 PAR_1_1_VDD075CPU 4.57849263885e-11
L_8_219 PAR_1_3_VDD075CPU n1267 3.31463180028e-06
R_8_219 n1267 PAR_1_1_VDD075CPU 242.640576171
G0_220 PAR_1_3_VDD075CPU PAR_2_1_VSS PAR_1_3_VDD075CPU PAR_2_1_VSS -1.4275317294
C0_220 PAR_1_3_VDD075CPU PAR_2_1_VSS 1.14757611772e-10
R_1_220 PAR_1_3_VDD075CPU n1268 1.24179051664
C_1_220 n1268 PAR_2_1_VSS 2.09636020787e-11
L_2_220 PAR_1_3_VDD075CPU n1269 8.22434191934e-11
R_2_220 n1269 PAR_2_1_VSS 1.08316769848
R_3_220 PAR_1_3_VDD075CPU n1270 2.18186300159
C_3_220 n1270 PAR_2_1_VSS 1.22037063942e-10
L_4_220 PAR_1_3_VDD075CPU n1271 1.16831174128e-09
R_4_220 n1271 PAR_2_1_VSS 2.34673219678
R_5_220 PAR_1_3_VDD075CPU n1272 6.6112638763
C_5_220 n1272 PAR_2_1_VSS 2.22668952269e-10
L_6_220 PAR_1_3_VDD075CPU n1273 5.41508600184e-08
R_6_220 n1273 PAR_2_1_VSS 12.7894916823
R_7_220 PAR_1_3_VDD075CPU n1274 78.9764771163
C_7_220 n1274 PAR_2_1_VSS 1.81003956179e-10
G0_221 PAR_1_3_VDD075CPU PAR_2_1_VDD075CPU PAR_1_3_VDD075CPU PAR_2_1_VDD075CPU -2.77362893107
C0_221 PAR_1_3_VDD075CPU PAR_2_1_VDD075CPU 9.68896162338e-11
R_1_221 PAR_1_3_VDD075CPU n1275 0.436866245356
C_1_221 n1275 PAR_2_1_VDD075CPU 5.6584149605e-11
L_2_221 PAR_1_3_VDD075CPU n1276 2.37445484859e-11
R_2_221 n1276 PAR_2_1_VDD075CPU 0.404525818923
R_3_221 PAR_1_3_VDD075CPU n1277 2.68238592853
C_3_221 n1277 PAR_2_1_VDD075CPU 4.5106710201e-11
L_4_221 PAR_1_3_VDD075CPU n1278 1.26138607633e-09
R_4_221 n1278 PAR_2_1_VDD075CPU 3.98264269991
R_5_221 PAR_1_3_VDD075CPU n1279 9.58803808595
C_5_221 n1279 PAR_2_1_VDD075CPU 9.11789630896e-11
L_6_221 PAR_1_3_VDD075CPU n1280 5.00157490907e-08
R_6_221 n1280 PAR_2_1_VDD075CPU 20.4332469786
R_7_221 PAR_1_3_VDD075CPU n1281 133.337940002
C_7_221 n1281 PAR_2_1_VDD075CPU 9.18794558702e-11
L_8_221 PAR_1_3_VDD075CPU n1282 0.000441271408254
R_8_221 n1282 PAR_2_1_VDD075CPU 633.008128784
G0_222 PAR_1_3_VDD075CPU PAR_0_2_VSS PAR_1_3_VDD075CPU PAR_0_2_VSS -0.229888573048
C0_222 PAR_1_3_VDD075CPU PAR_0_2_VSS 1.56785141387e-10
R_1_222 PAR_1_3_VDD075CPU n1283 0.116310084219
C_1_222 n1283 PAR_0_2_VSS 2.79796374344e-10
R_2_222 PAR_1_3_VDD075CPU n1284 1.08366513475
C_2_222 n1284 PAR_0_2_VSS 5.88180902315e-11
L_3_222 PAR_1_3_VDD075CPU n1285 1.86803646472e-09
R_3_222 n1285 PAR_0_2_VSS 4.6075940567
L_4_222 PAR_1_3_VDD075CPU n1286 1.97719899215e-07
R_4_222 n1286 PAR_0_2_VSS 77.7873097577
R_5_222 PAR_1_3_VDD075CPU n1287 29.7077566079
C_5_222 n1287 PAR_0_2_VSS 2.50404078764e-10
R0_223 PAR_1_3_VDD075CPU PAR_0_2_VDD075CPU 0.393186324355
C0_223 PAR_1_3_VDD075CPU PAR_0_2_VDD075CPU 1.46132748874e-10
L_1_223 PAR_1_3_VDD075CPU n1288 8.44817672378e-12
R_1_223 n1288 PAR_0_2_VDD075CPU 0.22351302258
L_2_223 PAR_1_3_VDD075CPU n1289 9.01495870317e-11
R_2_223 n1289 PAR_0_2_VDD075CPU 1.2126962109
L_3_223 PAR_1_3_VDD075CPU n1290 1.49589682049e-09
R_3_223 n1290 PAR_0_2_VDD075CPU 8.8984974188
L_4_223 PAR_1_3_VDD075CPU n1291 3.07212801891e-08
R_4_223 n1291 PAR_0_2_VDD075CPU 64.6452338128
L_5_223 PAR_1_3_VDD075CPU n1292 1.33449605725e-06
R_5_223 n1292 PAR_0_2_VDD075CPU 510.584668551
L_6_223 PAR_1_3_VDD075CPU n1293 0.000180210870759
R_6_223 n1293 PAR_0_2_VDD075CPU 3977.03284009
G0_224 PAR_1_3_VDD075CPU PAR_1_2_VSS PAR_1_3_VDD075CPU PAR_1_2_VSS -0.263290696223
C0_224 PAR_1_3_VDD075CPU PAR_1_2_VSS 1.21436890656e-10
R_1_224 PAR_1_3_VDD075CPU n1294 0.0271215412552
C_1_224 n1294 PAR_1_2_VSS 1.48032574684e-09
L_2_224 PAR_1_3_VDD075CPU n1295 3.7064698297e-10
R_2_224 n1295 PAR_1_2_VSS 3.90896596122
R_3_224 PAR_1_3_VDD075CPU n1296 77.5765260785
C_3_224 n1296 PAR_1_2_VSS 9.75100446602e-12
L_4_224 PAR_1_3_VDD075CPU n1297 1.28464362594e-06
R_4_224 n1297 PAR_1_2_VSS 133.894476531
R0_225 PAR_1_3_VDD075CPU PAR_1_2_VDD075CPU 0.00816258125167
C0_225 PAR_1_3_VDD075CPU PAR_1_2_VDD075CPU 8.7043621023e-11
L_1_225 PAR_1_3_VDD075CPU n1298 1.25736759207e-12
R_1_225 n1298 PAR_1_2_VDD075CPU 0.0583113922918
L_2_225 PAR_1_3_VDD075CPU n1299 6.54130533944e-13
R_2_225 n1299 PAR_1_2_VDD075CPU 0.0165087299293
L_3_225 PAR_1_3_VDD075CPU n1300 5.02327452706e-10
R_3_225 n1300 PAR_1_2_VDD075CPU 4.17191536395
L_4_225 PAR_1_3_VDD075CPU n1301 1.14181078849e-08
R_4_225 n1301 PAR_1_2_VDD075CPU 31.4731185895
L_5_225 PAR_1_3_VDD075CPU n1302 5.72776475135e-07
R_5_225 n1302 PAR_1_2_VDD075CPU 325.588525774
L_6_225 PAR_1_3_VDD075CPU n1303 9.92603997967e-05
R_6_225 n1303 PAR_1_2_VDD075CPU 4925.51795808
G0_226 PAR_1_3_VDD075CPU PAR_2_2_VSS PAR_1_3_VDD075CPU PAR_2_2_VSS -0.0374184717637
C0_226 PAR_1_3_VDD075CPU PAR_2_2_VSS 2.75858017318e-11
R_1_226 PAR_1_3_VDD075CPU n1304 0.187168877424
C_1_226 n1304 PAR_2_2_VSS 1.15103160107e-10
L_2_226 PAR_1_3_VDD075CPU n1305 2.36360161693e-08
R_2_226 n1305 PAR_2_2_VSS 111.376900584
L_3_226 PAR_1_3_VDD075CPU n1306 4.68863647039e-08
R_3_226 n1306 PAR_2_2_VSS 47.5421305704
L_4_226 PAR_1_3_VDD075CPU n1307 1.25632415382e-06
R_4_226 n1307 PAR_2_2_VSS 135.026085255
G0_227 PAR_1_3_VDD075CPU PAR_2_2_VDD075CPU PAR_1_3_VDD075CPU PAR_2_2_VDD075CPU -0.236380670577
C0_227 PAR_1_3_VDD075CPU PAR_2_2_VDD075CPU 1.72746754093e-11
R_1_227 PAR_1_3_VDD075CPU n1308 4.2304643504
C_1_227 n1308 PAR_2_2_VDD075CPU 4.80421793914e-12
L_2_227 PAR_1_3_VDD075CPU n1309 3.57000535168e-10
R_2_227 n1309 PAR_2_2_VDD075CPU 4.59162560944
L_3_227 PAR_1_3_VDD075CPU n1310 1.0602416379e-08
R_3_227 n1310 PAR_2_2_VDD075CPU 61.8672818169
L_4_227 PAR_1_3_VDD075CPU n1311 2.15728042726e-07
R_4_227 n1311 PAR_2_2_VDD075CPU 447.341348073
L_5_227 PAR_1_3_VDD075CPU n1312 1.78890715672e-05
R_5_227 n1312 PAR_2_2_VDD075CPU 5695.11071761
G0_228 PAR_1_3_VDD075CPU PAR_0_3_VSS PAR_1_3_VDD075CPU PAR_0_3_VSS -0.03112948025
C0_228 PAR_1_3_VDD075CPU PAR_0_3_VSS 1.89398037872e-10
R_1_228 PAR_1_3_VDD075CPU n1313 0.00862565939458
C_1_228 n1313 PAR_0_3_VSS 2.56512195566e-09
R_2_228 PAR_1_3_VDD075CPU n1314 0.0174866186031
C_2_228 n1314 PAR_0_3_VSS 2.41504679093e-09
R_3_228 PAR_1_3_VDD075CPU n1315 1.9882467211
C_3_228 n1315 PAR_0_3_VSS 7.79886563205e-11
L_4_228 PAR_1_3_VDD075CPU n1316 4.38929487849e-08
R_4_228 n1316 PAR_0_3_VSS 32.1238872372
R_5_228 PAR_1_3_VDD075CPU n1317 34.1442895831
C_5_228 n1317 PAR_0_3_VSS 2.51822402618e-10
R0_229 PAR_1_3_VDD075CPU PAR_0_3_VDD075CPU 0.00494720058231
C0_229 PAR_1_3_VDD075CPU PAR_0_3_VDD075CPU 4.14819886507e-11
L_1_229 PAR_1_3_VDD075CPU n1318 3.8471993067e-13
R_1_229 n1318 PAR_0_3_VDD075CPU 0.0168900839414
L_2_229 PAR_1_3_VDD075CPU n1319 8.35396696058e-13
R_2_229 n1319 PAR_0_3_VDD075CPU 0.0206761766957
L_3_229 PAR_1_3_VDD075CPU n1320 3.13903115039e-10
R_3_229 n1320 PAR_0_3_VDD075CPU 2.50676694137
L_4_229 PAR_1_3_VDD075CPU n1321 7.80018455358e-09
R_4_229 n1321 PAR_0_3_VDD075CPU 24.9880932571
L_5_229 PAR_1_3_VDD075CPU n1322 4.53865976114e-07
R_5_229 n1322 PAR_0_3_VDD075CPU 372.842019837
L_6_229 PAR_1_3_VDD075CPU n1323 1.39985286656e-05
R_6_229 n1323 PAR_0_3_VDD075CPU 1820.87855404
G0_230 PAR_1_3_VDD075CPU PAR_1_3_VSS PAR_1_3_VDD075CPU PAR_1_3_VSS -0.0319825071506
R_1_230 PAR_1_3_VDD075CPU n1324 0.000759917038625
C_1_230 n1324 PAR_1_3_VSS 2.36097191315e-08
R_2_230 PAR_1_3_VDD075CPU n1325 0.000636873758641
C_2_230 n1325 PAR_1_3_VSS 5.93842474675e-08
R_3_230 PAR_1_3_VDD075CPU n1326 0.178529750752
C_3_230 n1326 PAR_1_3_VSS 5.64595506606e-10
R_4_230 PAR_1_3_VDD075CPU n1327 0.642503674096
C_4_230 n1327 PAR_1_3_VSS 5.45795763748e-10
R_5_230 PAR_1_3_VDD075CPU n1328 4.67210636348
C_5_230 n1328 PAR_1_3_VSS 3.11393579858e-10
L_6_230 PAR_1_3_VDD075CPU n1329 3.33610082668e-07
R_6_230 n1329 PAR_1_3_VSS 31.2670895547
G0_231 PAR_1_3_VDD075CPU PAR_0_0_VSS PAR_1_3_VDD075CPU PAR_0_0_VSS -2.67367634653
C0_231 PAR_1_3_VDD075CPU PAR_0_0_VSS 2.29210548948e-10
R_1_231 PAR_1_3_VDD075CPU n1330 0.0206473420835
C_1_231 n1330 PAR_0_0_VSS 9.04376991514e-10
L_2_231 PAR_1_3_VDD075CPU n1331 4.29711076081e-11
R_2_231 n1331 PAR_0_0_VSS 0.474651414194
L_3_231 PAR_1_3_VDD075CPU n1332 5.68216420223e-10
R_3_231 n1332 PAR_0_0_VSS 1.76408198463
R_4_231 PAR_1_3_VDD075CPU n1333 20.3173875792
C_4_231 n1333 PAR_0_0_VSS 3.5610039915e-11
R_5_231 PAR_1_3_VDD075CPU n1334 214.37327046
C_5_231 n1334 PAR_0_0_VSS 7.6046097436e-11
.ENDS

