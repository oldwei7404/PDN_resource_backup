********************************************
* Ansys RedHawk-SC Chip Power Model [ Ver 2.00 ]
* Generated at Mar 08 11:59:16 2024
* Version: 2023 R1.2p1  RHEL7 (Mar 21 00:06:37 2023)
* Run directory:  /fs/mm_imp48/MM/PI/R0.7/RedHawk-SC/03_240203_wDFT_for_STAPI/MAMMOTH/v2023_R1.3_20230801/CPM_VDD075NNE_4x2_Flat/gp/asim_power_scratch.gv_rmv.240308033705.0j356unl
* CPM Options:
* perform powermodel -nx 4 -ny 2 -no_afs -noglobal_gnd -pincurrent -emi -plocnames
* Copyright (c) 2002-2023 ANSYS, Inc.
* Presimulation time  0.000000ps
********************************************


* Partitioning of flip chip bump pad area - Die Top View
* ------------------------------------
* | (0 Ny) | (1 Ny) | .... | (Nx Ny) |
* ------------------------------------
* | (0 ..) | (1 ..) | .... | (Nx ..) |
* ------------------------------------
* | (0  1) | (1  1) | .... | (Nx  1) |
* ------------------------------------
* | (0  0) | (1  0) | .... | (Nx  0) |
* ------------------------------------
* Begin Chip Package Protocol --->

.subckt adsPowerModel
+ PAR_0_0_VDD075NNE PAR_1_0_VSS PAR_1_0_VDD075NNE PAR_2_0_VSS PAR_2_0_VDD075NNE
+ PAR_3_0_VSS PAR_3_0_VDD075NNE PAR_0_1_VSS PAR_0_1_VDD075NNE PAR_1_1_VSS
+ PAR_1_1_VDD075NNE PAR_2_1_VSS PAR_2_1_VDD075NNE PAR_3_1_VSS PAR_3_1_VDD075NNE
+ PAR_0_0_VSS

* Xpdn
* + PAR_0_0_VDD075NNE PAR_1_0_VSS PAR_1_0_VDD075NNE PAR_2_0_VSS PAR_2_0_VDD075NNE
* + PAR_3_0_VSS PAR_3_0_VDD075NNE PAR_0_1_VSS PAR_0_1_VDD075NNE PAR_1_1_VSS
* + PAR_1_1_VDD075NNE PAR_2_1_VSS PAR_2_1_VDD075NNE PAR_3_1_VSS PAR_3_1_VDD075NNE
* + PAR_0_0_VSS
* + PowerModel

* CPM Port Name | Average current (A) | Max. magnitude of current | Net voltage *
* PAR_0_0_VSS -3.73536 5.10844 0
* PAR_0_0_VDD075NNE 4.17578 7.74687 0.7125
* PAR_1_0_VSS -3.80984 5.35321 0
* PAR_1_0_VDD075NNE 3.79172 6.90731 0.7125
* PAR_2_0_VSS -3.69164 5.30191 0
* PAR_2_0_VDD075NNE 4.07567 7.36738 0.7125
* PAR_3_0_VSS -5.05814 8.04883 0
* PAR_3_0_VDD075NNE 5.31282 11.5551 0.7125
* PAR_0_1_VSS -19.6666 27.8128 0
* PAR_0_1_VDD075NNE 21.8669 38.7293 0.7125
* PAR_1_1_VSS -19.8214 30.4777 0
* PAR_1_1_VDD075NNE 19.75 36.6949 0.7125
* PAR_2_1_VSS -18.9626 27.6987 0
* PAR_2_1_VDD075NNE 22.0788 40.0233 0.7125
* PAR_3_1_VSS -19.1364 26.4486 0
* PAR_3_1_VDD075NNE 19.8665 33.9918 0.7125
* Average power = 71.9042 W.

* .SUBCKT PowerModel PAR_0_0_VDD075NNE PAR_1_0_VSS PAR_1_0_VDD075NNE PAR_2_0_VSS PAR_2_0_VDD075NNE
* + PAR_3_0_VSS PAR_3_0_VDD075NNE PAR_0_1_VSS PAR_0_1_VDD075NNE PAR_1_1_VSS
* + PAR_1_1_VDD075NNE PAR_2_1_VSS PAR_2_1_VDD075NNE PAR_3_1_VSS PAR_3_1_VDD075NNE
* + PAR_0_0_VSS
**********************************************************
* Ansys RedHawk-SC Chip Power Model [Accurate RC reduction]
* Model Subcircuit of Die PDN
* Copyright (c) 2002-2023 ANSYS, Inc.
**********************************************************

* No connection to global ground (Spice node 0) *
G0_1 PAR_0_0_VDD075NNE PAR_0_0_VSS PAR_0_0_VDD075NNE PAR_0_0_VSS -0.0184733093274
C0_1 PAR_0_0_VDD075NNE PAR_0_0_VSS 1.76518976662e-09
R_1_1 PAR_0_0_VDD075NNE n17 0.00023783977852
C_1_1 n17 PAR_0_0_VSS 5.93229268207e-08
R_2_1 PAR_0_0_VDD075NNE n18 0.000567318472783
C_2_1 n18 PAR_0_0_VSS 5.53865144867e-08
R_3_1 PAR_0_0_VDD075NNE n19 0.164732465067
C_3_1 n19 PAR_0_0_VSS 5.91605095037e-10
R_4_1 PAR_0_0_VDD075NNE n20 1.26295098032
R_7_1 PAR_0_0_VDD075NNE n20 1778000
C_4_1 n20 PAR_0_0_VSS 2.83672626402e-10
R_5_1 PAR_0_0_VDD075NNE n21 7.01645410484
R_8_1 PAR_0_0_VDD075NNE n21 1889000
C_5_1 n21 PAR_0_0_VSS 2.73268520813e-10
L_6_1 PAR_0_0_VDD075NNE n22 6.25714680802e-07
R_6_1 n22 PAR_0_0_VSS 54.1321445097
G0_2 PAR_1_0_VSS PAR_0_0_VDD075NNE PAR_1_0_VSS PAR_0_0_VDD075NNE -0.0558402389441
C0_2 PAR_1_0_VSS PAR_0_0_VDD075NNE 2.04397933727e-10
R_1_2 PAR_1_0_VSS n23 0.00440445437612
C_1_2 n23 PAR_0_0_VDD075NNE 3.20434372253e-09
R_2_2 PAR_1_0_VSS n24 0.0085152105941
C_2_2 n24 PAR_0_0_VDD075NNE 3.61256432818e-09
L_3_2 PAR_1_0_VSS n25 4.94108732509e-09
R_3_2 n25 PAR_0_0_VDD075NNE 24.7700425165
R_4_2 PAR_1_0_VSS n26 5.8466521971
R_9_2 PAR_1_0_VSS n26 1666000
C_4_2 n26 PAR_0_0_VDD075NNE 7.09382995646e-11
R_5_2 PAR_1_0_VSS n27 11.0735572606
R_10_2 PAR_1_0_VSS n27 1484000
C_5_2 n27 PAR_0_0_VDD075NNE 1.62207588336e-10
L_6_2 PAR_1_0_VSS n28 6.8552676963e-07
R_6_2 n28 PAR_0_0_VDD075NNE 64.645860991
R0_3 PAR_1_0_VSS PAR_0_0_VSS 0.00291787960813
L_1_3 PAR_1_0_VSS n29 1.42356097241e-13
R_1_3 n29 PAR_0_0_VSS 0.00596202697554
R_2_3 PAR_1_0_VSS n30 0.292414042655
C_2_3 n30 PAR_0_0_VSS 6.80099356271e-10
L_3_3 PAR_1_0_VSS n31 7.05642405359e-11
R_3_3 n31 PAR_0_0_VSS 0.181821965604
L_4_3 PAR_1_0_VSS n32 5.69297052758e-10
R_4_3 n32 PAR_0_0_VSS 0.161727071201
L_5_3 PAR_1_0_VSS n33 4.15267569018e-09
R_5_3 n33 PAR_0_0_VSS 0.421878738207
R0_4 PAR_1_0_VDD075NNE PAR_0_0_VDD075NNE 0.00344995455113
C0_4 PAR_1_0_VDD075NNE PAR_0_0_VDD075NNE 7.02017726412e-11
L_1_4 PAR_1_0_VDD075NNE n34 1.25873189806e-13
R_1_4 n34 PAR_0_0_VDD075NNE 0.00767694841026
L_2_4 PAR_1_0_VDD075NNE n35 4.3160027081e-13
R_2_4 n35 PAR_0_0_VDD075NNE 0.0134719580126
L_3_4 PAR_1_0_VDD075NNE n36 3.49462309769e-10
R_3_4 n36 PAR_0_0_VDD075NNE 3.98515797627
L_4_4 PAR_1_0_VDD075NNE n37 2.10535081218e-08
R_4_4 n37 PAR_0_0_VDD075NNE 57.7169286788
L_5_4 PAR_1_0_VDD075NNE n38 1.94837732047e-07
R_5_4 n38 PAR_0_0_VDD075NNE 157.736248977
L_6_4 PAR_1_0_VDD075NNE n39 4.93694304289e-05
R_6_4 n39 PAR_0_0_VDD075NNE 3633.16227217
G0_5 PAR_1_0_VDD075NNE PAR_1_0_VSS PAR_1_0_VDD075NNE PAR_1_0_VSS -0.013535635826
C0_5 PAR_1_0_VDD075NNE PAR_1_0_VSS 1.20459420361e-09
R_1_5 PAR_1_0_VDD075NNE n40 0.00023786896752
C_1_5 n40 PAR_1_0_VSS 5.53751034899e-08
R_2_5 PAR_1_0_VDD075NNE n41 0.000579957361358
C_2_5 n41 PAR_1_0_VSS 5.14861723937e-08
R_3_5 PAR_1_0_VDD075NNE n42 0.0916047212506
C_3_5 n42 PAR_1_0_VSS 7.88264476134e-10
R_4_5 PAR_1_0_VDD075NNE n43 2.97517254599
C_4_5 n43 PAR_1_0_VSS 1.17053469256e-10
R_5_5 PAR_1_0_VDD075NNE n44 9.36796986655
C_5_5 n44 PAR_1_0_VSS 1.66206326686e-10
L_6_5 PAR_1_0_VDD075NNE n45 8.22345041192e-07
R_6_5 n45 PAR_1_0_VSS 73.8790379495
G0_6 PAR_1_0_VDD075NNE PAR_0_0_VSS PAR_1_0_VDD075NNE PAR_0_0_VSS -0.0690790583589
C0_6 PAR_1_0_VDD075NNE PAR_0_0_VSS 1.26693911951e-10
R_1_6 PAR_1_0_VDD075NNE n46 0.0145612037667
C_1_6 n46 PAR_0_0_VSS 1.18949538638e-09
R_2_6 PAR_1_0_VDD075NNE n47 0.0211248790038
C_2_6 n47 PAR_0_0_VSS 1.53165524197e-09
L_3_6 PAR_1_0_VDD075NNE n48 2.44363040324e-09
R_3_6 n48 PAR_0_0_VSS 21.6614888507
R_4_6 PAR_1_0_VDD075NNE n49 5.48560002656
C_4_6 n49 PAR_0_0_VSS 7.33820126332e-11
R_5_6 PAR_1_0_VDD075NNE n50 12.2527426783
C_5_6 n50 PAR_0_0_VSS 1.77265419077e-10
L_6_6 PAR_1_0_VDD075NNE n51 4.25901408535e-07
R_6_6 n51 PAR_0_0_VSS 43.641093837
G0_7 PAR_2_0_VSS PAR_0_0_VDD075NNE PAR_2_0_VSS PAR_0_0_VDD075NNE -1.73636010747
C0_7 PAR_2_0_VSS PAR_0_0_VDD075NNE 1.29029114606e-10
R_1_7 PAR_2_0_VSS n52 0.787071331393
C_1_7 n52 PAR_0_0_VDD075NNE 1.75764123692e-11
L_2_7 PAR_2_0_VSS n53 2.35299644743e-11
R_2_7 n53 PAR_0_0_VDD075NNE 0.657513268774
R_3_7 PAR_2_0_VSS n54 5.38070605778
C_3_7 n54 PAR_0_0_VDD075NNE 2.83124322631e-11
L_4_7 PAR_2_0_VSS n55 4.5681822521e-09
R_4_7 n55 PAR_0_0_VDD075NNE 12.0308331141
R_5_7 PAR_2_0_VSS n56 4.44054635892
C_5_7 n56 PAR_0_0_VDD075NNE 1.71950700151e-10
L_6_7 PAR_2_0_VSS n57 1.21163817619e-08
R_6_7 n57 PAR_0_0_VDD075NNE 8.84119842145
R_7_7 PAR_2_0_VSS n58 18.2546692466
C_7_7 n58 PAR_0_0_VDD075NNE 1.64110626043e-10
L_8_7 PAR_2_0_VSS n59 4.79180818014e-07
R_8_7 n59 PAR_0_0_VDD075NNE 51.9435894597
R0_8 PAR_2_0_VSS PAR_1_0_VSS 0.00331887189638
L_1_8 PAR_2_0_VSS n60 1.19366202074e-13
R_1_8 n60 PAR_1_0_VSS 0.00514797718304
L_2_8 PAR_2_0_VSS n61 1.7098014768e-11
R_2_8 n61 PAR_1_0_VSS 0.20921456864
L_3_8 PAR_2_0_VSS n62 7.58148868207e-11
R_3_8 n62 PAR_1_0_VSS 0.244200709222
L_4_8 PAR_2_0_VSS n63 3.92674291374e-10
R_4_8 n63 PAR_1_0_VSS 0.583666572048
L_5_8 PAR_2_0_VSS n64 5.71140127114e-10
R_5_8 n64 PAR_1_0_VSS 0.257301210297
L_6_8 PAR_2_0_VSS n65 7.70123447147e-09
R_6_8 n65 PAR_1_0_VSS 0.885580342424
G0_9 PAR_2_0_VSS PAR_1_0_VDD075NNE PAR_2_0_VSS PAR_1_0_VDD075NNE -0.00852747614327
C0_9 PAR_2_0_VSS PAR_1_0_VDD075NNE 1.05794858591e-10
R_1_9 PAR_2_0_VSS n66 0.0116218625806
C_1_9 n66 PAR_1_0_VDD075NNE 1.77418466795e-09
R_2_9 PAR_2_0_VSS n67 0.0515358902426
C_2_9 n67 PAR_1_0_VDD075NNE 7.44719357351e-10
R_3_9 PAR_2_0_VSS n68 7.32163409851
C_3_9 n68 PAR_1_0_VDD075NNE 1.92358159315e-11
R_4_9 PAR_2_0_VSS n69 7.73677060224
C_4_9 n69 PAR_1_0_VDD075NNE 5.59246370885e-11
R_5_9 PAR_2_0_VSS n70 20.5994483472
C_5_9 n70 PAR_1_0_VDD075NNE 7.92715362294e-11
L_6_9 PAR_2_0_VSS n71 1.17378400151e-06
R_6_9 n71 PAR_1_0_VDD075NNE 117.267949379
R0_10 PAR_2_0_VSS PAR_0_0_VSS 0.901489099116
C0_10 PAR_2_0_VSS PAR_0_0_VSS 1.71355160611e-10
R_1_10 PAR_2_0_VSS n72 0.805030512053
C_1_10 n72 PAR_0_0_VSS 7.41427551296e-11
R_2_10 PAR_2_0_VSS n73 1.48785630196
C_2_10 n73 PAR_0_0_VSS 3.38450170223e-10
R_3_10 PAR_2_0_VSS n74 0.449635433249
C_3_10 n74 PAR_0_0_VSS 4.06416834943e-09
L_4_10 PAR_2_0_VSS n75 5.23173290892e-09
R_4_10 n75 PAR_0_0_VSS 1.04925710734
L_5_10 PAR_2_0_VSS n76 8.11861892065e-09
R_5_10 n76 PAR_0_0_VSS 0.841582601229
G0_11 PAR_2_0_VDD075NNE PAR_0_0_VDD075NNE PAR_2_0_VDD075NNE PAR_0_0_VDD075NNE -5.60200154636
C0_11 PAR_2_0_VDD075NNE PAR_0_0_VDD075NNE 1.107653288e-10
R_1_11 PAR_2_0_VDD075NNE n77 0.223158024302
C_1_11 n77 PAR_0_0_VDD075NNE 5.8816999555e-11
L_2_11 PAR_2_0_VDD075NNE n78 7.06894987052e-12
R_2_11 n78 PAR_0_0_VDD075NNE 0.193425625416
R_3_11 PAR_2_0_VDD075NNE n79 1.04051303389
C_3_11 n79 PAR_0_0_VDD075NNE 7.04054177582e-11
L_4_11 PAR_2_0_VDD075NNE n80 5.00321703597e-10
R_4_11 n80 PAR_0_0_VDD075NNE 2.97412848038
R_5_11 PAR_2_0_VDD075NNE n81 7.97991922576
C_5_11 n81 PAR_0_0_VDD075NNE 5.07512695272e-11
L_6_11 PAR_2_0_VDD075NNE n82 1.05013319745e-08
R_6_11 n82 PAR_0_0_VDD075NNE 11.0398636423
R_7_11 PAR_2_0_VDD075NNE n83 28.9912599153
C_7_11 n83 PAR_0_0_VDD075NNE 6.42453994404e-11
L_8_11 PAR_2_0_VDD075NNE n84 1.74247169236e-06
R_8_11 n84 PAR_0_0_VDD075NNE 193.762701377
G0_12 PAR_2_0_VDD075NNE PAR_1_0_VSS PAR_2_0_VDD075NNE PAR_1_0_VSS -0.0172654845886
C0_12 PAR_2_0_VDD075NNE PAR_1_0_VSS 2.10265965687e-10
R_1_12 PAR_2_0_VDD075NNE n85 0.00351009807921
C_1_12 n85 PAR_1_0_VSS 4.50510198974e-09
R_2_12 PAR_2_0_VDD075NNE n86 0.0131319102368
C_2_12 n86 PAR_1_0_VSS 2.5947969669e-09
R_3_12 PAR_2_0_VDD075NNE n87 2.4601780125
C_3_12 n87 PAR_1_0_VSS 4.12049228341e-11
R_4_12 PAR_2_0_VDD075NNE n88 5.93292498323
C_4_12 n88 PAR_1_0_VSS 7.04087381315e-11
R_5_12 PAR_2_0_VDD075NNE n89 10.7371160082
C_5_12 n89 PAR_1_0_VSS 1.59850543378e-10
L_6_12 PAR_2_0_VDD075NNE n90 5.82822533047e-07
R_6_12 n90 PAR_1_0_VSS 57.9190106655
R0_13 PAR_2_0_VDD075NNE PAR_1_0_VDD075NNE 0.00372480345999
C0_13 PAR_2_0_VDD075NNE PAR_1_0_VDD075NNE 6.95098514495e-11
L_1_13 PAR_2_0_VDD075NNE n91 9.70342160209e-14
R_1_13 n91 PAR_1_0_VDD075NNE 0.00595976323333
L_2_13 PAR_2_0_VDD075NNE n92 6.97519372043e-13
R_2_13 n92 PAR_1_0_VDD075NNE 0.0204058415365
L_3_13 PAR_2_0_VDD075NNE n93 1.63473101459e-10
R_3_13 n93 PAR_1_0_VDD075NNE 1.9593092863
L_4_13 PAR_2_0_VDD075NNE n94 2.55532879083e-08
R_4_13 n94 PAR_1_0_VDD075NNE 62.2560346305
L_5_13 PAR_2_0_VDD075NNE n95 3.01032673146e-07
R_5_13 n95 PAR_1_0_VDD075NNE 202.351072505
L_6_13 PAR_2_0_VDD075NNE n96 0.00505428670637
R_6_13 n96 PAR_1_0_VDD075NNE 2514.27858737
G0_14 PAR_2_0_VDD075NNE PAR_2_0_VSS PAR_2_0_VDD075NNE PAR_2_0_VSS -0.00822230689573
C0_14 PAR_2_0_VDD075NNE PAR_2_0_VSS 1.01336490872e-09
R_1_14 PAR_2_0_VDD075NNE n97 0.000244325490111
C_1_14 n97 PAR_2_0_VSS 5.19040840923e-08
R_2_14 PAR_2_0_VDD075NNE n98 0.000539886254275
C_2_14 n98 PAR_2_0_VSS 5.39284374003e-08
R_3_14 PAR_2_0_VDD075NNE n99 0.0545565491407
C_3_14 n99 PAR_2_0_VSS 1.10638742617e-09
R_4_14 PAR_2_0_VDD075NNE n100 4.58656043468
C_4_14 n100 PAR_2_0_VSS 8.1835775903e-11
R_5_14 PAR_2_0_VDD075NNE n101 15.5379305227
C_5_14 n101 PAR_2_0_VSS 9.19617248285e-11
L_6_14 PAR_2_0_VDD075NNE n102 1.3330386604e-06
R_6_14 n102 PAR_2_0_VSS 121.620319112
G0_15 PAR_2_0_VDD075NNE PAR_0_0_VSS PAR_2_0_VDD075NNE PAR_0_0_VSS -0.0259597126108
C0_15 PAR_2_0_VDD075NNE PAR_0_0_VSS 1.68340341558e-10
R_1_15 PAR_2_0_VDD075NNE n103 0.403107860473
C_1_15 n103 PAR_0_0_VSS 7.38860184016e-11
R_2_15 PAR_2_0_VDD075NNE n104 6.2635479708
C_2_15 n104 PAR_0_0_VSS 6.24134802987e-11
R_3_15 PAR_2_0_VDD075NNE n105 12.6005039709
C_3_15 n105 PAR_0_0_VSS 1.69907956876e-10
L_4_15 PAR_2_0_VDD075NNE n106 3.69582274918e-07
R_4_15 n106 PAR_0_0_VSS 38.5212229977
G0_16 PAR_3_0_VSS PAR_0_0_VDD075NNE PAR_3_0_VSS PAR_0_0_VDD075NNE -1.03087844606
C0_16 PAR_3_0_VSS PAR_0_0_VDD075NNE 2.47765365155e-10
R_1_16 PAR_3_0_VSS n107 0.0386551015824
C_1_16 n107 PAR_0_0_VDD075NNE 4.91504112891e-10
R_2_16 PAR_3_0_VSS n108 0.25326248063
C_2_16 n108 PAR_0_0_VDD075NNE 1.94920964382e-10
L_3_16 PAR_3_0_VSS n109 1.18696150457e-10
R_3_16 n109 PAR_0_0_VDD075NNE 0.970046468207
R_4_16 PAR_3_0_VSS n110 3.34919894431
C_4_16 n110 PAR_0_0_VDD075NNE 1.2032536471e-10
R_5_16 PAR_3_0_VSS n111 3.59130791768
C_5_16 n111 PAR_0_0_VDD075NNE 2.64312033408e-10
R_6_16 PAR_3_0_VSS n112 37.1760145234
C_6_16 n112 PAR_0_0_VDD075NNE 3.03583386347e-10
R0_17 PAR_3_0_VSS PAR_1_0_VSS 0.144667054321
C0_17 PAR_3_0_VSS PAR_1_0_VSS 2.48879199003e-10
R_1_17 PAR_3_0_VSS n113 0.0882435225141
C_1_17 n113 PAR_1_0_VSS 2.90578886522e-10
R_2_17 PAR_3_0_VSS n114 0.0982780379293
C_2_17 n114 PAR_1_0_VSS 9.80591767247e-10
R_3_17 PAR_3_0_VSS n115 0.46591920642
C_3_17 n115 PAR_1_0_VSS 6.3015103023e-10
R_4_17 PAR_3_0_VSS n116 0.4142244423
C_4_17 n116 PAR_1_0_VSS 1.81963415004e-09
R_5_17 PAR_3_0_VSS n117 0.193466099465
C_5_17 n117 PAR_1_0_VSS 1.89042040059e-08
R_6_17 PAR_3_0_VSS n118 0.403170676022
C_6_17 n118 PAR_1_0_VSS 2.5156857764e-08
G0_18 PAR_3_0_VSS PAR_1_0_VDD075NNE PAR_3_0_VSS PAR_1_0_VDD075NNE -0.546927021078
C0_18 PAR_3_0_VSS PAR_1_0_VDD075NNE 2.11815479442e-10
R_1_18 PAR_3_0_VSS n119 0.0465460971028
C_1_18 n119 PAR_1_0_VDD075NNE 3.40732187603e-10
R_2_18 PAR_3_0_VSS n120 0.235807052646
C_2_18 n120 PAR_1_0_VDD075NNE 2.00136899221e-10
L_3_18 PAR_3_0_VSS n121 2.27734372506e-10
R_3_18 n121 PAR_1_0_VDD075NNE 1.82839748852
R_4_18 PAR_3_0_VSS n122 3.12339367557
C_4_18 n122 PAR_1_0_VDD075NNE 1.39967371027e-10
R_5_18 PAR_3_0_VSS n123 4.39745800775
C_5_18 n123 PAR_1_0_VDD075NNE 2.34190148745e-10
R_6_18 PAR_3_0_VSS n124 33.7179624832
C_6_18 n124 PAR_1_0_VDD075NNE 2.97875148654e-10
R0_19 PAR_3_0_VSS PAR_2_0_VSS 0.00271375136643
L_1_19 PAR_3_0_VSS n125 1.63456971188e-13
R_1_19 n125 PAR_2_0_VSS 0.00667984748722
R_2_19 PAR_3_0_VSS n126 0.292087358214
C_2_19 n126 PAR_2_0_VSS 6.20626104683e-10
L_3_19 PAR_3_0_VSS n127 8.83573767794e-11
R_3_19 n127 PAR_2_0_VSS 0.222368260463
L_4_19 PAR_3_0_VSS n128 9.39903633912e-10
R_4_19 n128 PAR_2_0_VSS 0.574227868333
R_5_19 PAR_3_0_VSS n129 0.842590082739
C_5_19 n129 PAR_2_0_VSS 8.92370066471e-09
R_6_19 PAR_3_0_VSS n130 2.62136232093
C_6_19 n130 PAR_2_0_VSS 5.45402563217e-09
C0_20 PAR_3_0_VSS PAR_2_0_VDD075NNE 1.55245636237e-10
R_1_20 PAR_3_0_VSS n131 0.00402820562117
C_1_20 n131 PAR_2_0_VDD075NNE 3.2307516007e-09
R_2_20 PAR_3_0_VSS n132 0.00767951140059
C_2_20 n132 PAR_2_0_VDD075NNE 4.04265875791e-09
R_3_20 PAR_3_0_VSS n133 2.00522681014
C_3_20 n133 PAR_2_0_VDD075NNE 3.17536923741e-10
R_4_20 PAR_3_0_VSS n134 14.9306361473
C_4_20 n134 PAR_2_0_VDD075NNE 1.24393980206e-10
R_5_20 PAR_3_0_VSS n135 32.931965856
C_5_20 n135 PAR_2_0_VDD075NNE 3.17133217182e-10
R0_21 PAR_3_0_VSS PAR_0_0_VSS 1.1289722211
C0_21 PAR_3_0_VSS PAR_0_0_VSS 2.05162536744e-10
R_1_21 PAR_3_0_VSS n136 0.0981909960091
C_1_21 n136 PAR_0_0_VSS 6.11884231533e-10
R_2_21 PAR_3_0_VSS n137 0.0780110346836
C_2_21 n137 PAR_0_0_VSS 1.62472025923e-09
R_3_21 PAR_3_0_VSS n138 0.137907036574
C_3_21 n138 PAR_0_0_VSS 4.18914304872e-09
L_4_21 PAR_3_0_VSS n139 4.69019912345e-10
R_4_21 n139 PAR_0_0_VSS 0.519579587893
R_5_21 PAR_3_0_VSS n140 0.0699233414118
C_5_21 n140 PAR_0_0_VSS 4.58229324382e-08
R_6_21 PAR_3_0_VSS n141 0.250184728397
C_6_21 n141 PAR_0_0_VSS 3.95189675836e-08
G0_22 PAR_3_0_VDD075NNE PAR_0_0_VDD075NNE PAR_3_0_VDD075NNE PAR_0_0_VDD075NNE -6.00322865031
C0_22 PAR_3_0_VDD075NNE PAR_0_0_VDD075NNE 1.93231366157e-10
R_1_22 PAR_3_0_VDD075NNE n142 0.0607231899624
C_1_22 n142 PAR_0_0_VDD075NNE 1.00020822726e-10
L_2_22 PAR_3_0_VDD075NNE n143 7.77938379916e-12
R_2_22 n143 PAR_0_0_VDD075NNE 0.23810267162
L_3_22 PAR_3_0_VDD075NNE n144 3.66169646996e-11
R_3_22 n144 PAR_0_0_VDD075NNE 0.59060250699
L_4_22 PAR_3_0_VDD075NNE n145 3.34367541742e-09
R_4_22 n145 PAR_0_0_VDD075NNE 17.5737149396
L_5_22 PAR_3_0_VDD075NNE n146 1.12214946209e-08
R_5_22 n146 PAR_0_0_VDD075NNE 24.7973067311
L_6_22 PAR_3_0_VDD075NNE n147 1.00823699588e-07
R_6_22 n147 PAR_0_0_VDD075NNE 81.2831805347
L_7_22 PAR_3_0_VDD075NNE n148 7.76165387484e-06
R_7_22 n148 PAR_0_0_VDD075NNE 1426.22926879
G0_23 PAR_3_0_VDD075NNE PAR_1_0_VSS PAR_3_0_VDD075NNE PAR_1_0_VSS -0.00706653928367
C0_23 PAR_3_0_VDD075NNE PAR_1_0_VSS 2.31843563465e-10
R_1_23 PAR_3_0_VDD075NNE n149 0.124444384032
C_1_23 n149 PAR_1_0_VSS 1.69885473773e-10
R_2_23 PAR_3_0_VDD075NNE n150 3.68366668514
C_2_23 n150 PAR_1_0_VSS 1.40947745013e-10
L_3_23 PAR_3_0_VDD075NNE n151 6.90278290905e-06
R_3_23 n151 PAR_1_0_VSS 141.511908851
G0_24 PAR_3_0_VDD075NNE PAR_1_0_VDD075NNE PAR_3_0_VDD075NNE PAR_1_0_VDD075NNE -39.5797884622
C0_24 PAR_3_0_VDD075NNE PAR_1_0_VDD075NNE 1.49817120621e-10
R_1_24 PAR_3_0_VDD075NNE n152 0.0309177804883
C_1_24 n152 PAR_1_0_VDD075NNE 1.51431738723e-09
L_2_24 PAR_3_0_VDD075NNE n153 1.45605087947e-12
R_2_24 n153 PAR_1_0_VDD075NNE 0.026224862211
R_3_24 PAR_3_0_VDD075NNE n154 0.152695118815
C_3_24 n154 PAR_1_0_VDD075NNE 6.21910191828e-10
L_4_24 PAR_3_0_VDD075NNE n155 2.46347000263e-10
R_4_24 n155 PAR_1_0_VDD075NNE 0.839673889751
R_5_24 PAR_3_0_VDD075NNE n156 1.52406157083
C_5_24 n156 PAR_1_0_VDD075NNE 4.14107737483e-10
L_6_24 PAR_3_0_VDD075NNE n157 6.07026303662e-09
R_6_24 n157 PAR_1_0_VDD075NNE 3.96414228391
R_7_24 PAR_3_0_VDD075NNE n158 32.4665474427
C_7_24 n158 PAR_1_0_VDD075NNE 2.34211485382e-10
L_8_24 PAR_3_0_VDD075NNE n159 0.00114456087245
R_8_24 n159 PAR_1_0_VDD075NNE 204.683916338
G0_25 PAR_3_0_VDD075NNE PAR_2_0_VSS PAR_3_0_VDD075NNE PAR_2_0_VSS -0.0117413168942
C0_25 PAR_3_0_VDD075NNE PAR_2_0_VSS 1.63971815882e-10
R_1_25 PAR_3_0_VDD075NNE n160 0.015690637882
C_1_25 n160 PAR_2_0_VSS 1.04192653819e-09
R_2_25 PAR_3_0_VDD075NNE n161 0.0203285705968
C_2_25 n161 PAR_2_0_VSS 1.55502482786e-09
R_3_25 PAR_3_0_VDD075NNE n162 4.33251633348
C_3_25 n162 PAR_2_0_VSS 2.64043769885e-11
R_4_25 PAR_3_0_VDD075NNE n163 6.45492206113
C_4_25 n163 PAR_2_0_VSS 6.7461224899e-11
R_5_25 PAR_3_0_VDD075NNE n164 8.33160079777
C_5_25 n164 PAR_2_0_VSS 2.51074365244e-10
L_6_25 PAR_3_0_VDD075NNE n165 7.74558305466e-07
R_6_25 n165 PAR_2_0_VSS 85.1692968532
R0_26 PAR_3_0_VDD075NNE PAR_2_0_VDD075NNE 0.00369397455833
C0_26 PAR_3_0_VDD075NNE PAR_2_0_VDD075NNE 1.03260814407e-10
L_1_26 PAR_3_0_VDD075NNE n166 1.32421591374e-13
R_1_26 n166 PAR_2_0_VDD075NNE 0.00737142976822
L_2_26 PAR_3_0_VDD075NNE n167 5.63097197505e-13
R_2_26 n167 PAR_2_0_VDD075NNE 0.0166433089866
L_3_26 PAR_3_0_VDD075NNE n168 1.61529181816e-10
R_3_26 n168 PAR_2_0_VDD075NNE 1.80781348627
L_4_26 PAR_3_0_VDD075NNE n169 7.10381339237e-09
R_4_26 n169 PAR_2_0_VDD075NNE 19.9643935072
L_5_26 PAR_3_0_VDD075NNE n170 6.0221315203e-08
R_5_26 n170 PAR_2_0_VDD075NNE 58.0912644973
L_6_26 PAR_3_0_VDD075NNE n171 4.38196895002e-06
R_6_26 n171 PAR_2_0_VDD075NNE 1013.74814283
C0_27 PAR_3_0_VDD075NNE PAR_3_0_VSS 3.02644468619e-09
R_1_27 PAR_3_0_VDD075NNE n172 0.000204761246726
C_1_27 n172 PAR_3_0_VSS 7.93831287206e-08
R_2_27 PAR_3_0_VDD075NNE n173 0.000718219799106
C_2_27 n173 PAR_3_0_VSS 5.20120676543e-08
R_3_27 PAR_3_0_VDD075NNE n174 0.0739095005333
C_3_27 n174 PAR_3_0_VSS 1.75470549411e-09
R_4_27 PAR_3_0_VDD075NNE n175 0.105676729785
C_4_27 n175 PAR_3_0_VSS 3.00619188224e-09
R_5_27 PAR_3_0_VDD075NNE n176 0.662755581137
C_5_27 n176 PAR_3_0_VSS 1.51061624733e-09
R_6_27 PAR_3_0_VDD075NNE n177 4.69106973945
C_6_27 n177 PAR_3_0_VSS 1.14542411332e-09
G0_28 PAR_3_0_VDD075NNE PAR_0_0_VSS PAR_3_0_VDD075NNE PAR_0_0_VSS -0.049110519817
C0_28 PAR_3_0_VDD075NNE PAR_0_0_VSS 2.32597499794e-10
R_1_28 PAR_3_0_VDD075NNE n178 0.0801077118254
C_1_28 n178 PAR_0_0_VSS 3.66662409802e-10
R_2_28 PAR_3_0_VDD075NNE n179 2.93290464068
C_2_28 n179 PAR_0_0_VSS 1.45621951981e-10
L_3_28 PAR_3_0_VDD075NNE n180 1.18030551847e-07
R_3_28 n180 PAR_0_0_VSS 20.3622347661
G0_29 PAR_0_1_VSS PAR_0_0_VDD075NNE PAR_0_1_VSS PAR_0_0_VDD075NNE -0.533381970171
C0_29 PAR_0_1_VSS PAR_0_0_VDD075NNE 2.24738945944e-10
R_1_29 PAR_0_1_VSS n181 0.0274966551905
C_1_29 n181 PAR_0_0_VDD075NNE 8.78413673117e-10
R_2_29 PAR_0_1_VSS n182 0.10073260673
C_2_29 n182 PAR_0_0_VDD075NNE 4.66651947696e-10
L_3_29 PAR_0_1_VSS n183 8.32612716698e-10
R_3_29 n183 PAR_0_0_VDD075NNE 2.56939928512
L_4_29 PAR_0_1_VSS n184 7.12304621127e-09
R_4_29 n184 PAR_0_0_VDD075NNE 7.49352942527
L_5_29 PAR_0_1_VSS n185 3.92921498277e-07
R_5_29 n185 PAR_0_0_VDD075NNE 93.1317310987
R0_30 PAR_0_1_VSS PAR_1_0_VSS 0.152800586609
C0_30 PAR_0_1_VSS PAR_1_0_VSS 2.4119203537e-10
R_1_30 PAR_0_1_VSS n186 0.588714751349
C_1_30 n186 PAR_1_0_VSS 7.63393703029e-11
R_2_30 PAR_0_1_VSS n187 0.274628461196
C_2_30 n187 PAR_1_0_VSS 5.02200127863e-10
R_3_30 PAR_0_1_VSS n188 0.270013107752
C_3_30 n188 PAR_1_0_VSS 1.29999838279e-09
R_4_30 PAR_0_1_VSS n189 1.58381352968
C_4_30 n189 PAR_1_0_VSS 5.91967687644e-10
R_5_30 PAR_0_1_VSS n190 1.11471002326
C_5_30 n190 PAR_1_0_VSS 1.76354596514e-09
L_6_30 PAR_0_1_VSS n191 3.67205494803e-08
R_6_30 n191 PAR_1_0_VSS 3.88731161546
G0_31 PAR_0_1_VSS PAR_1_0_VDD075NNE PAR_0_1_VSS PAR_1_0_VDD075NNE -0.417738739382
C0_31 PAR_0_1_VSS PAR_1_0_VDD075NNE 2.05700214866e-10
R_1_31 PAR_0_1_VSS n192 0.247691148687
C_1_31 n192 PAR_1_0_VDD075NNE 9.5640617953e-11
R_2_31 PAR_0_1_VSS n193 3.92306565768
C_2_31 n193 PAR_1_0_VDD075NNE 2.12733365149e-11
L_3_31 PAR_0_1_VSS n194 1.28508291156e-09
R_3_31 n194 PAR_1_0_VDD075NNE 4.11319687422
L_4_31 PAR_0_1_VSS n195 5.3257763722e-09
R_4_31 n195 PAR_1_0_VDD075NNE 8.25806030328
L_5_31 PAR_0_1_VSS n196 2.92690096926e-08
R_5_31 n196 PAR_1_0_VDD075NNE 19.8572863497
L_6_31 PAR_0_1_VSS n197 2.65466362892e-06
R_6_31 n197 PAR_1_0_VDD075NNE 315.887312952
G0_32 PAR_0_1_VSS PAR_2_0_VSS PAR_0_1_VSS PAR_2_0_VSS -0.139187709397
C0_32 PAR_0_1_VSS PAR_2_0_VSS 2.0909871394e-10
R_1_32 PAR_0_1_VSS n198 0.626665150414
C_1_32 n198 PAR_2_0_VSS 4.71387550774e-11
R_2_32 PAR_0_1_VSS n199 0.907730790795
C_2_32 n199 PAR_2_0_VSS 1.66186263036e-10
R_3_32 PAR_0_1_VSS n200 0.365654479872
C_3_32 n200 PAR_2_0_VSS 1.0405313558e-09
R_4_32 PAR_0_1_VSS n201 2.32211452496
C_4_32 n201 PAR_2_0_VSS 4.06124319849e-10
R_5_32 PAR_0_1_VSS n202 2.31921427747
C_5_32 n202 PAR_2_0_VSS 8.08471345658e-10
L_6_32 PAR_0_1_VSS n203 6.75320713057e-08
R_6_32 n203 PAR_2_0_VSS 7.1845357843
G0_33 PAR_0_1_VSS PAR_2_0_VDD075NNE PAR_0_1_VSS PAR_2_0_VDD075NNE -0.429728099619
C0_33 PAR_0_1_VSS PAR_2_0_VDD075NNE 2.12697782205e-10
R_1_33 PAR_0_1_VSS n204 0.382034888517
C_1_33 n204 PAR_2_0_VDD075NNE 6.1140000625e-11
R_2_33 PAR_0_1_VSS n205 3.46384541192
C_2_33 n205 PAR_2_0_VDD075NNE 2.80809536507e-11
L_3_33 PAR_0_1_VSS n206 1.30982442368e-09
R_3_33 n206 PAR_2_0_VDD075NNE 4.13346680902
L_4_33 PAR_0_1_VSS n207 4.92505246303e-09
R_4_33 n207 PAR_2_0_VDD075NNE 7.71192943792
L_5_33 PAR_0_1_VSS n208 2.66010479439e-08
R_5_33 n208 PAR_2_0_VDD075NNE 18.2900151233
L_6_33 PAR_0_1_VSS n209 2.43364930071e-06
R_6_33 n209 PAR_2_0_VDD075NNE 289.305358294
R0_34 PAR_0_1_VSS PAR_3_0_VSS 83509.3238527
C0_34 PAR_0_1_VSS PAR_3_0_VSS 2.85184964107e-10
R_1_34 PAR_0_1_VSS n210 0.0716061532028
C_1_34 n210 PAR_3_0_VSS 5.87246050645e-10
R_2_34 PAR_0_1_VSS n211 0.0471117583716
C_2_34 n211 PAR_3_0_VSS 2.63361701995e-09
R_3_34 PAR_0_1_VSS n212 0.0697287881817
C_3_34 n212 PAR_3_0_VSS 3.61975441247e-09
R_4_34 PAR_0_1_VSS n213 0.148078313756
C_4_34 n213 PAR_3_0_VSS 3.48916624222e-09
R_5_34 PAR_0_1_VSS n214 0.328530447091
C_5_34 n214 PAR_3_0_VSS 3.42783493598e-09
R_6_34 PAR_0_1_VSS n215 2.20632466602
C_6_34 n215 PAR_3_0_VSS 4.43513080649e-09
G0_35 PAR_0_1_VSS PAR_3_0_VDD075NNE PAR_0_1_VSS PAR_3_0_VDD075NNE -1.24439317985
C0_35 PAR_0_1_VSS PAR_3_0_VDD075NNE 2.6952875632e-10
R_1_35 PAR_0_1_VSS n216 0.0618020119338
C_1_35 n216 PAR_3_0_VDD075NNE 2.84127033646e-10
R_2_35 PAR_0_1_VSS n217 0.251217178634
C_2_35 n217 PAR_3_0_VDD075NNE 1.84037562376e-10
L_3_35 PAR_0_1_VSS n218 4.80295885401e-10
R_3_35 n218 PAR_3_0_VDD075NNE 1.44019739435
L_4_35 PAR_0_1_VSS n219 1.40820317386e-09
R_4_35 n219 PAR_3_0_VDD075NNE 2.35893175895
L_5_35 PAR_0_1_VSS n220 1.19691772034e-08
R_5_35 n220 PAR_3_0_VDD075NNE 8.27352638422
L_6_35 PAR_0_1_VSS n221 1.40624169062e-06
R_6_35 n221 PAR_3_0_VDD075NNE 190.266867193
R0_36 PAR_0_1_VSS PAR_0_0_VSS 0.00825483243315
C0_36 PAR_0_1_VSS PAR_0_0_VSS 1.56907532394e-10
L_1_36 PAR_0_1_VSS n222 3.51158094893e-13
R_1_36 n222 PAR_0_0_VSS 0.0153623504424
L_2_36 PAR_0_1_VSS n223 3.48176184702e-12
R_2_36 n223 PAR_0_0_VSS 0.0777718669476
R_3_36 PAR_0_1_VSS n224 0.153162645413
C_3_36 n224 PAR_0_0_VSS 1.06327983191e-09
R_4_36 PAR_0_1_VSS n225 0.184466174847
C_4_36 n225 PAR_0_0_VSS 1.98885442745e-09
R_5_36 PAR_0_1_VSS n226 0.851504245225
C_5_36 n226 PAR_0_0_VSS 2.43020237604e-09
L_6_36 PAR_0_1_VSS n227 2.81639422228e-08
R_6_36 n227 PAR_0_0_VSS 2.91267624339
R0_37 PAR_0_1_VDD075NNE PAR_0_0_VDD075NNE 0.00774451837393
C0_37 PAR_0_1_VDD075NNE PAR_0_0_VDD075NNE 2.04711946647e-10
L_1_37 PAR_0_1_VDD075NNE n228 2.80147832888e-13
R_1_37 n228 PAR_0_0_VDD075NNE 0.0133817409811
L_2_37 PAR_0_1_VDD075NNE n229 1.37404117869e-12
R_2_37 n229 PAR_0_0_VDD075NNE 0.0337911414401
L_3_37 PAR_0_1_VDD075NNE n230 1.79858384436e-10
R_3_37 n230 PAR_0_0_VDD075NNE 1.99948107905
L_4_37 PAR_0_1_VDD075NNE n231 3.83425373235e-08
R_4_37 n231 PAR_0_0_VDD075NNE 70.9660791043
L_5_37 PAR_0_1_VDD075NNE n232 3.74663985914e-07
R_5_37 n232 PAR_0_0_VDD075NNE 208.748189424
L_6_37 PAR_0_1_VDD075NNE n233 0.00398388324455
R_6_37 n233 PAR_0_0_VDD075NNE 2356.82718441
G0_38 PAR_0_1_VDD075NNE PAR_1_0_VSS PAR_0_1_VDD075NNE PAR_1_0_VSS -0.348331820071
C0_38 PAR_0_1_VDD075NNE PAR_1_0_VSS 2.48421742758e-10
R_1_38 PAR_0_1_VDD075NNE n234 0.089964321464
C_1_38 n234 PAR_1_0_VSS 2.03016962351e-10
R_2_38 PAR_0_1_VDD075NNE n235 0.324599439048
C_2_38 n235 PAR_1_0_VSS 1.32238244585e-10
L_3_38 PAR_0_1_VDD075NNE n236 4.0528103131e-10
R_3_38 n236 PAR_1_0_VSS 3.09026434392
R_4_38 PAR_0_1_VDD075NNE n237 9.95565193571
C_4_38 n237 PAR_1_0_VSS 4.72271074747e-11
R_5_38 PAR_0_1_VDD075NNE n238 9.44688308122
C_5_38 n238 PAR_1_0_VSS 1.85185415471e-10
L_6_38 PAR_0_1_VDD075NNE n239 3.95587894048e-07
R_6_38 n239 PAR_1_0_VSS 40.4286865129
G0_39 PAR_0_1_VDD075NNE PAR_1_0_VDD075NNE PAR_0_1_VDD075NNE PAR_1_0_VDD075NNE -0.279947989014
C0_39 PAR_0_1_VDD075NNE PAR_1_0_VDD075NNE 1.65508110361e-10
L_1_39 PAR_0_1_VDD075NNE n240 4.98174341418e-12
R_1_39 n240 PAR_1_0_VDD075NNE 0.216353342919
L_2_39 PAR_0_1_VDD075NNE n241 1.57203305154e-11
R_2_39 n241 PAR_1_0_VDD075NNE 0.296125277978
R_3_39 PAR_0_1_VDD075NNE n242 3.79562674615
C_3_39 n242 PAR_1_0_VDD075NNE 3.81404694962e-11
L_4_39 PAR_0_1_VDD075NNE n243 7.81371036594e-09
R_4_39 n243 PAR_1_0_VDD075NNE 11.4235305811
R_5_39 PAR_0_1_VDD075NNE n244 60.654258995
C_5_39 n244 PAR_1_0_VDD075NNE 3.81444581215e-11
G0_40 PAR_0_1_VDD075NNE PAR_2_0_VSS PAR_0_1_VDD075NNE PAR_2_0_VSS -2.77133719841
C0_40 PAR_0_1_VDD075NNE PAR_2_0_VSS 1.73903414268e-10
R_1_40 PAR_0_1_VDD075NNE n245 0.404981002651
C_1_40 n245 PAR_2_0_VSS 3.93817941071e-11
L_2_40 PAR_0_1_VDD075NNE n246 1.16910725114e-11
R_2_40 n246 PAR_2_0_VSS 0.367341258785
R_3_40 PAR_0_1_VDD075NNE n247 6.43358777333
C_3_40 n247 PAR_2_0_VSS 1.89415036626e-11
R_4_40 PAR_0_1_VDD075NNE n248 66.9086544919
C_4_40 n248 PAR_2_0_VSS 6.14525010366e-12
R_5_40 PAR_0_1_VDD075NNE n249 7.59269423247
C_5_40 n249 PAR_2_0_VSS 1.74232116991e-10
L_6_40 PAR_0_1_VDD075NNE n250 6.03883063555e-08
R_6_40 n250 PAR_2_0_VSS 24.5170232958
L_7_40 PAR_0_1_VDD075NNE n251 1.11503871952e-06
R_7_40 n251 PAR_2_0_VSS 120.701488657
G0_41 PAR_0_1_VDD075NNE PAR_2_0_VDD075NNE PAR_0_1_VDD075NNE PAR_2_0_VDD075NNE -8.41986311652
C0_41 PAR_0_1_VDD075NNE PAR_2_0_VDD075NNE 1.44135172502e-10
R_1_41 PAR_0_1_VDD075NNE n252 0.155224632036
C_1_41 n252 PAR_2_0_VDD075NNE 9.95633685572e-11
L_2_41 PAR_0_1_VDD075NNE n253 5.05639852042e-12
R_2_41 n253 PAR_2_0_VDD075NNE 0.132361054552
R_3_41 PAR_0_1_VDD075NNE n254 0.590264925054
C_3_41 n254 PAR_2_0_VDD075NNE 1.36367588436e-10
L_4_41 PAR_0_1_VDD075NNE n255 2.25618245086e-10
R_4_41 n255 PAR_2_0_VDD075NNE 1.43809297293
R_5_41 PAR_0_1_VDD075NNE n256 4.54951020475
C_5_41 n256 PAR_2_0_VDD075NNE 9.22574711824e-11
L_6_41 PAR_0_1_VDD075NNE n257 5.96062155281e-09
R_6_41 n257 PAR_2_0_VDD075NNE 6.22904015179
R_7_41 PAR_0_1_VDD075NNE n258 15.7163032263
C_7_41 n258 PAR_2_0_VDD075NNE 1.17244283924e-10
L_8_41 PAR_0_1_VDD075NNE n259 1.04699792333e-06
R_8_41 n259 PAR_2_0_VDD075NNE 115.386386656
G0_42 PAR_0_1_VDD075NNE PAR_3_0_VSS PAR_0_1_VDD075NNE PAR_3_0_VSS -2.05136177052
C0_42 PAR_0_1_VDD075NNE PAR_3_0_VSS 3.0811417201e-10
R_1_42 PAR_0_1_VDD075NNE n260 0.0259560775931
C_1_42 n260 PAR_3_0_VSS 6.62211704642e-10
R_2_42 PAR_0_1_VDD075NNE n261 0.152543329185
C_2_42 n261 PAR_3_0_VSS 3.29444822083e-10
L_3_42 PAR_0_1_VDD075NNE n262 6.91689706545e-11
R_3_42 n262 PAR_3_0_VSS 0.487481053617
R_4_42 PAR_0_1_VDD075NNE n263 2.92688941773
C_4_42 n263 PAR_3_0_VSS 1.80357775963e-10
R_5_42 PAR_0_1_VDD075NNE n264 3.89261735184
C_5_42 n264 PAR_3_0_VSS 2.87318205766e-10
R_6_42 PAR_0_1_VDD075NNE n265 21.556059608
C_6_42 n265 PAR_3_0_VSS 4.52900345199e-10
G0_43 PAR_0_1_VDD075NNE PAR_3_0_VDD075NNE PAR_0_1_VDD075NNE PAR_3_0_VDD075NNE -8.13291799721
C0_43 PAR_0_1_VDD075NNE PAR_3_0_VDD075NNE 2.11301502887e-10
R_1_43 PAR_0_1_VDD075NNE n266 0.0222301710961
C_1_43 n266 PAR_3_0_VDD075NNE 1.82211899257e-10
L_2_43 PAR_0_1_VDD075NNE n267 5.56395609962e-12
R_2_43 n267 PAR_3_0_VDD075NNE 0.163513332608
L_3_43 PAR_0_1_VDD075NNE n268 3.59684238963e-11
R_3_43 n268 PAR_3_0_VDD075NNE 0.521085612348
L_4_43 PAR_0_1_VDD075NNE n269 3.87498270894e-09
R_4_43 n269 PAR_3_0_VDD075NNE 20.6231331214
L_5_43 PAR_0_1_VDD075NNE n270 1.40642110062e-08
R_5_43 n270 PAR_3_0_VDD075NNE 28.5941495188
L_6_43 PAR_0_1_VDD075NNE n271 9.21041590123e-08
R_6_43 n271 PAR_3_0_VDD075NNE 72.3615210171
L_7_43 PAR_0_1_VDD075NNE n272 6.00681025603e-06
R_7_43 n272 PAR_3_0_VDD075NNE 1058.39530327
G0_44 PAR_0_1_VDD075NNE PAR_0_1_VSS PAR_0_1_VDD075NNE PAR_0_1_VSS -0.192826358099
C0_44 PAR_0_1_VDD075NNE PAR_0_1_VSS 8.53076969449e-10
R_1_44 PAR_0_1_VDD075NNE n273 0.000416532984881
C_1_44 n273 PAR_0_1_VSS 3.16760686876e-08
R_2_44 PAR_0_1_VDD075NNE n274 0.000250174102863
C_2_44 n274 PAR_0_1_VSS 1.32413451779e-07
R_3_44 PAR_0_1_VDD075NNE n275 0.00226571825166
C_3_44 n275 PAR_0_1_VSS 2.17010908422e-08
R_4_44 PAR_0_1_VDD075NNE n276 0.142959811992
C_4_44 n276 PAR_0_1_VSS 1.06899154396e-09
L_5_44 PAR_0_1_VDD075NNE n277 4.91743509898e-09
R_5_44 n277 PAR_0_1_VSS 5.68857459434
L_6_44 PAR_0_1_VDD075NNE n278 2.18410437276e-07
R_6_44 n278 PAR_0_1_VSS 58.7012908365
G0_45 PAR_0_1_VDD075NNE PAR_0_0_VSS PAR_0_1_VDD075NNE PAR_0_0_VSS -0.0237441160563
C0_45 PAR_0_1_VDD075NNE PAR_0_0_VSS 2.30151267713e-10
R_1_45 PAR_0_1_VDD075NNE n279 0.00645262753473
C_1_45 n279 PAR_0_0_VSS 2.3590304234e-09
R_2_45 PAR_0_1_VDD075NNE n280 0.0143316234433
C_2_45 n280 PAR_0_0_VSS 2.6155030439e-09
R_3_45 PAR_0_1_VDD075NNE n281 7.15990037115
C_3_45 n281 PAR_0_0_VSS 1.99008130153e-10
L_4_45 PAR_0_1_VDD075NNE n282 5.19515739273e-07
R_4_45 n282 PAR_0_0_VSS 42.1156907653
G0_46 PAR_1_1_VSS PAR_0_0_VDD075NNE PAR_1_1_VSS PAR_0_0_VDD075NNE -0.639440985573
C0_46 PAR_1_1_VSS PAR_0_0_VDD075NNE 2.44930699299e-10
R_1_46 PAR_1_1_VSS n283 0.114362209545
C_1_46 n283 PAR_0_0_VDD075NNE 1.69352188264e-10
R_2_46 PAR_1_1_VSS n284 0.837071987633
C_2_46 n284 PAR_0_0_VDD075NNE 7.73358767736e-11
L_3_46 PAR_1_1_VSS n285 8.511774279e-10
R_3_46 n285 PAR_0_0_VDD075NNE 2.8196090167
L_4_46 PAR_1_1_VSS n286 2.89385118725e-09
R_4_46 n286 PAR_0_0_VDD075NNE 4.91282824488
L_5_46 PAR_1_1_VSS n287 1.881432597e-08
R_5_46 n287 PAR_0_0_VDD075NNE 13.0390364502
L_6_46 PAR_1_1_VSS n288 1.78953236925e-06
R_6_46 n288 PAR_0_0_VDD075NNE 220.246657696
R0_47 PAR_1_1_VSS PAR_1_0_VSS 0.00866772135584
C0_47 PAR_1_1_VSS PAR_1_0_VSS 1.31343871679e-10
L_1_47 PAR_1_1_VSS n289 4.1399737724e-13
R_1_47 n289 PAR_1_0_VSS 0.0151373425282
R_2_47 PAR_1_1_VSS n290 0.214014492132
C_2_47 n290 PAR_1_0_VSS 8.7551678651e-10
R_3_47 PAR_1_1_VSS n291 0.260835587633
C_3_47 n291 PAR_1_0_VSS 1.65245214855e-09
R_4_47 PAR_1_1_VSS n292 0.683541171631
C_4_47 n292 PAR_1_0_VSS 2.56736146728e-09
L_5_47 PAR_1_1_VSS n293 3.19562993602e-08
R_5_47 n293 PAR_1_0_VSS 3.27792264526
G0_48 PAR_1_1_VSS PAR_1_0_VDD075NNE PAR_1_1_VSS PAR_1_0_VDD075NNE -0.457202297276
C0_48 PAR_1_1_VSS PAR_1_0_VDD075NNE 2.14950601225e-10
R_1_48 PAR_1_1_VSS n294 0.0302843047442
C_1_48 n294 PAR_1_0_VDD075NNE 8.14353680817e-10
R_2_48 PAR_1_1_VSS n295 0.204336165065
C_2_48 n295 PAR_1_0_VDD075NNE 2.77524296904e-10
L_3_48 PAR_1_1_VSS n296 1.19007764554e-09
R_3_48 n296 PAR_1_0_VDD075NNE 2.95832599936
L_4_48 PAR_1_1_VSS n297 1.02441283992e-08
R_4_48 n297 PAR_1_0_VDD075NNE 8.87007587877
L_5_48 PAR_1_1_VSS n298 9.46201394288e-07
R_5_48 n298 PAR_1_0_VDD075NNE 155.407721282
R0_49 PAR_1_1_VSS PAR_2_0_VSS 0.204931888383
C0_49 PAR_1_1_VSS PAR_2_0_VSS 2.24107571487e-10
L_1_49 PAR_1_1_VSS n299 2.43291873477e-11
R_1_49 n299 PAR_2_0_VSS 0.618407148082
R_2_49 PAR_1_1_VSS n300 0.791881774288
C_2_49 n300 PAR_2_0_VSS 1.93198421449e-10
R_3_49 PAR_1_1_VSS n301 0.27856278457
C_3_49 n301 PAR_2_0_VSS 1.40177349424e-09
R_4_49 PAR_1_1_VSS n302 1.59742044504
C_4_49 n302 PAR_2_0_VSS 7.13357842828e-10
R_5_49 PAR_1_1_VSS n303 2.67141007907
C_5_49 n303 PAR_2_0_VSS 7.80344708762e-10
L_6_49 PAR_1_1_VSS n304 5.25881865545e-08
R_6_49 n304 PAR_2_0_VSS 5.64771550482
G0_50 PAR_1_1_VSS PAR_2_0_VDD075NNE PAR_1_1_VSS PAR_2_0_VDD075NNE -0.471644215821
C0_50 PAR_1_1_VSS PAR_2_0_VDD075NNE 2.27783243545e-10
R_1_50 PAR_1_1_VSS n305 0.181503682481
C_1_50 n305 PAR_2_0_VDD075NNE 1.29924179742e-10
R_2_50 PAR_1_1_VSS n306 0.885324274925
C_2_50 n306 PAR_2_0_VDD075NNE 8.70561936707e-11
L_3_50 PAR_1_1_VSS n307 1.20112765707e-09
R_3_50 n307 PAR_2_0_VDD075NNE 2.96520869686
L_4_50 PAR_1_1_VSS n308 8.8658647721e-09
R_4_50 n308 PAR_2_0_VDD075NNE 8.30893674272
L_5_50 PAR_1_1_VSS n309 2.43854665537e-07
R_5_50 n309 PAR_2_0_VDD075NNE 88.4158119003
L_6_50 PAR_1_1_VSS n310 3.87095478128e-06
R_6_50 n310 PAR_2_0_VDD075NNE 365.32447784
R0_51 PAR_1_1_VSS PAR_3_0_VSS 75177.2931405
C0_51 PAR_1_1_VSS PAR_3_0_VSS 2.77915181416e-10
R_1_51 PAR_1_1_VSS n311 0.0827439678436
C_1_51 n311 PAR_3_0_VSS 3.5524256544e-10
R_2_51 PAR_1_1_VSS n312 0.0355942760825
C_2_51 n312 PAR_3_0_VSS 3.71560407835e-09
R_3_51 PAR_1_1_VSS n313 0.0541647451769
C_3_51 n313 PAR_3_0_VSS 5.33460472259e-09
R_4_51 PAR_1_1_VSS n314 0.146433790972
C_4_51 n314 PAR_3_0_VSS 4.09655119633e-09
R_5_51 PAR_1_1_VSS n315 0.317151624367
C_5_51 n315 PAR_3_0_VSS 3.73026179647e-09
R_6_51 PAR_1_1_VSS n316 1.78057972402
C_6_51 n316 PAR_3_0_VSS 5.52106890602e-09
G0_52 PAR_1_1_VSS PAR_3_0_VDD075NNE PAR_1_1_VSS PAR_3_0_VDD075NNE -1.42847486096
C0_52 PAR_1_1_VSS PAR_3_0_VDD075NNE 2.80858823144e-10
R_1_52 PAR_1_1_VSS n317 0.0499267143113
C_1_52 n317 PAR_3_0_VDD075NNE 3.42877110551e-10
R_2_52 PAR_1_1_VSS n318 0.216865692593
C_2_52 n318 PAR_3_0_VDD075NNE 2.80037857302e-10
L_3_52 PAR_1_1_VSS n319 3.79350642688e-10
R_3_52 n319 PAR_3_0_VDD075NNE 0.930900076799
L_4_52 PAR_1_1_VSS n320 3.14429136486e-09
R_4_52 n320 PAR_3_0_VDD075NNE 3.51908454535
L_5_52 PAR_1_1_VSS n321 2.88070744207e-08
R_5_52 n321 PAR_3_0_VDD075NNE 15.2428721257
L_6_52 PAR_1_1_VSS n322 2.02871359096e-06
R_6_52 n322 PAR_3_0_VDD075NNE 223.390476754
R0_53 PAR_1_1_VSS PAR_0_1_VSS 0.00243187871218
L_1_53 PAR_1_1_VSS n323 1.82955449737e-13
R_1_53 n323 PAR_0_1_VSS 0.00524640610369
R_2_53 PAR_1_1_VSS n324 0.0281420844981
C_2_53 n324 PAR_0_1_VSS 5.92331769677e-09
L_3_53 PAR_1_1_VSS n325 7.7620162967e-12
R_3_53 n325 PAR_0_1_VSS 0.0290397249635
L_4_53 PAR_1_1_VSS n326 2.99997173114e-10
R_4_53 n326 PAR_0_1_VSS 0.341770570067
L_5_53 PAR_1_1_VSS n327 2.27697872444e-08
R_5_53 n327 PAR_0_1_VSS 5.27741805686
G0_54 PAR_1_1_VSS PAR_0_1_VDD075NNE PAR_1_1_VSS PAR_0_1_VDD075NNE -1.04456080414
C0_54 PAR_1_1_VSS PAR_0_1_VDD075NNE 4.31219670883e-10
R_1_54 PAR_1_1_VSS n328 0.00554439278238
C_1_54 n328 PAR_0_1_VDD075NNE 3.83741482434e-09
R_2_54 PAR_1_1_VSS n329 0.00507874933162
C_2_54 n329 PAR_0_1_VDD075NNE 7.71689324641e-09
L_3_54 PAR_1_1_VSS n330 2.05085484084e-10
R_3_54 n330 PAR_0_1_VDD075NNE 1.26725827207
L_4_54 PAR_1_1_VSS n331 3.61371702118e-09
R_4_54 n331 PAR_0_1_VDD075NNE 4.29439398617
L_5_54 PAR_1_1_VSS n332 1.59104234949e-07
R_5_54 n332 PAR_0_1_VDD075NNE 44.2596271249
R0_55 PAR_1_1_VSS PAR_0_0_VSS 0.159464780128
C0_55 PAR_1_1_VSS PAR_0_0_VSS 2.3057702093e-10
R_1_55 PAR_1_1_VSS n333 0.36133922657
C_1_55 n333 PAR_0_0_VSS 9.48974366723e-11
R_2_55 PAR_1_1_VSS n334 0.151842900279
C_2_55 n334 PAR_0_0_VSS 8.81497255605e-10
R_3_55 PAR_1_1_VSS n335 0.178406563718
C_3_55 n335 PAR_0_0_VSS 1.49982552762e-09
R_4_55 PAR_1_1_VSS n336 0.244616603042
C_4_55 n336 PAR_0_0_VSS 1.70420222287e-09
R_5_55 PAR_1_1_VSS n337 0.692016956409
C_5_55 n337 PAR_0_0_VSS 3.06605524814e-09
L_6_55 PAR_1_1_VSS n338 2.16355402086e-08
R_6_55 n338 PAR_0_0_VSS 2.27337486085
G0_56 PAR_1_1_VDD075NNE PAR_0_0_VDD075NNE PAR_1_1_VDD075NNE PAR_0_0_VDD075NNE -0.246684077222
C0_56 PAR_1_1_VDD075NNE PAR_0_0_VDD075NNE 1.71491315317e-10
L_1_56 PAR_1_1_VDD075NNE n339 4.90592424562e-12
R_1_56 n339 PAR_0_0_VDD075NNE 0.199264377994
L_2_56 PAR_1_1_VDD075NNE n340 1.84256337621e-11
R_2_56 n340 PAR_0_0_VDD075NNE 0.335585014242
R_3_56 PAR_1_1_VDD075NNE n341 4.38651643171
C_3_56 n341 PAR_0_0_VDD075NNE 3.89763130067e-11
L_4_56 PAR_1_1_VDD075NNE n342 7.06639749495e-09
R_4_56 n342 PAR_0_0_VDD075NNE 10.1415404584
R_5_56 PAR_1_1_VDD075NNE n343 53.4395175023
C_5_56 n343 PAR_0_0_VDD075NNE 4.44073192226e-11
G0_57 PAR_1_1_VDD075NNE PAR_1_0_VSS PAR_1_1_VDD075NNE PAR_1_0_VSS -0.0254649386428
C0_57 PAR_1_1_VDD075NNE PAR_1_0_VSS 2.63685771055e-10
R_1_57 PAR_1_1_VDD075NNE n344 0.00621566918241
C_1_57 n344 PAR_1_0_VSS 2.70622317362e-09
R_2_57 PAR_1_1_VDD075NNE n345 0.0222995314062
C_2_57 n345 PAR_1_0_VSS 1.77527954932e-09
R_3_57 PAR_1_1_VDD075NNE n346 10.9422101094
C_3_57 n346 PAR_1_0_VSS 5.72311103075e-11
R_4_57 PAR_1_1_VDD075NNE n347 12.4749634669
C_4_57 n347 PAR_1_0_VSS 1.63844453772e-10
L_5_57 PAR_1_1_VDD075NNE n348 3.53625179672e-07
R_5_57 n348 PAR_1_0_VSS 39.269675284
R0_58 PAR_1_1_VDD075NNE PAR_1_0_VDD075NNE 0.00889067253361
C0_58 PAR_1_1_VDD075NNE PAR_1_0_VDD075NNE 1.57755847252e-10
L_1_58 PAR_1_1_VDD075NNE n349 2.75836795705e-13
R_1_58 n349 PAR_1_0_VDD075NNE 0.0136589431083
L_2_58 PAR_1_1_VDD075NNE n350 1.94160438672e-12
R_2_58 n350 PAR_1_0_VDD075NNE 0.0475770214894
L_3_58 PAR_1_1_VDD075NNE n351 4.17247837138e-10
R_3_58 n351 PAR_1_0_VDD075NNE 4.0744631999
L_4_58 PAR_1_1_VDD075NNE n352 3.99078576045e-08
R_4_58 n352 PAR_1_0_VDD075NNE 79.7199090148
L_5_58 PAR_1_1_VDD075NNE n353 4.03743453718e-07
R_5_58 n353 PAR_1_0_VDD075NNE 234.887122156
L_6_58 PAR_1_1_VDD075NNE n354 0.00762611031432
R_6_58 n354 PAR_1_0_VDD075NNE 1432.66562806
G0_59 PAR_1_1_VDD075NNE PAR_2_0_VSS PAR_1_1_VDD075NNE PAR_2_0_VSS -0.0116029322875
C0_59 PAR_1_1_VDD075NNE PAR_2_0_VSS 1.77640482186e-10
R_1_59 PAR_1_1_VDD075NNE n355 0.646759587205
C_1_59 n355 PAR_2_0_VSS 6.4327591362e-11
R_2_59 PAR_1_1_VDD075NNE n356 10.3463167253
C_2_59 n356 PAR_2_0_VSS 3.98319132945e-11
R_3_59 PAR_1_1_VDD075NNE n357 18.3020142647
C_3_59 n357 PAR_2_0_VSS 8.36740393578e-11
L_4_59 PAR_1_1_VDD075NNE n358 8.62136139765e-07
R_4_59 n358 PAR_2_0_VSS 86.1850881468
G0_60 PAR_1_1_VDD075NNE PAR_2_0_VDD075NNE PAR_1_1_VDD075NNE PAR_2_0_VDD075NNE -0.213635064332
C0_60 PAR_1_1_VDD075NNE PAR_2_0_VDD075NNE 1.46980400884e-10
L_1_60 PAR_1_1_VDD075NNE n359 4.06788668974e-12
R_1_60 n359 PAR_2_0_VDD075NNE 0.196205670147
L_2_60 PAR_1_1_VDD075NNE n360 1.81699679452e-11
R_2_60 n360 PAR_2_0_VDD075NNE 0.345082765193
R_3_60 PAR_1_1_VDD075NNE n361 5.04150955513
C_3_60 n361 PAR_2_0_VDD075NNE 3.09288652671e-11
L_4_60 PAR_1_1_VDD075NNE n362 7.80622422854e-09
R_4_60 n362 PAR_2_0_VDD075NNE 11.7590139395
R_5_60 PAR_1_1_VDD075NNE n363 65.4374217053
C_5_60 n363 PAR_2_0_VDD075NNE 3.43304243687e-11
G0_61 PAR_1_1_VDD075NNE PAR_3_0_VSS PAR_1_1_VDD075NNE PAR_3_0_VSS -1.28738967479
C0_61 PAR_1_1_VDD075NNE PAR_3_0_VSS 2.65202438664e-10
R_1_61 PAR_1_1_VDD075NNE n364 0.029036436112
C_1_61 n364 PAR_3_0_VSS 5.39036756146e-10
R_2_61 PAR_1_1_VDD075NNE n365 0.173317914994
C_2_61 n365 PAR_3_0_VSS 2.78730452647e-10
L_3_61 PAR_1_1_VDD075NNE n366 1.09923796447e-10
R_3_61 n366 PAR_3_0_VSS 0.776765587108
R_4_61 PAR_1_1_VDD075NNE n367 3.22503665211
C_4_61 n367 PAR_3_0_VSS 1.68147543366e-10
R_5_61 PAR_1_1_VDD075NNE n368 4.45794903246
C_5_61 n368 PAR_3_0_VSS 2.53444958981e-10
R_6_61 PAR_1_1_VDD075NNE n369 24.0922269101
C_6_61 n369 PAR_3_0_VSS 4.05809977084e-10
G0_62 PAR_1_1_VDD075NNE PAR_3_0_VDD075NNE PAR_1_1_VDD075NNE PAR_3_0_VDD075NNE -7.61145324669
C0_62 PAR_1_1_VDD075NNE PAR_3_0_VDD075NNE 1.71522726923e-10
R_1_62 PAR_1_1_VDD075NNE n370 0.0202774230105
C_1_62 n370 PAR_3_0_VDD075NNE 1.73607041266e-10
L_2_62 PAR_1_1_VDD075NNE n371 5.45336554951e-12
R_2_62 n371 PAR_3_0_VDD075NNE 0.183379888838
L_3_62 PAR_1_1_VDD075NNE n372 3.13301834979e-11
R_3_62 n372 PAR_3_0_VDD075NNE 0.497199924409
L_4_62 PAR_1_1_VDD075NNE n373 1.68307094881e-09
R_4_62 n373 PAR_3_0_VDD075NNE 11.8082474319
L_5_62 PAR_1_1_VDD075NNE n374 9.30728724164e-09
R_5_62 n374 PAR_3_0_VDD075NNE 27.8486597881
L_6_62 PAR_1_1_VDD075NNE n375 3.82537401388e-08
R_6_62 n375 PAR_3_0_VDD075NNE 51.6313360967
L_7_62 PAR_1_1_VDD075NNE n376 2.4624299126e-07
R_7_62 n376 PAR_3_0_VDD075NNE 149.879769503
L_8_62 PAR_1_1_VDD075NNE n377 2.08117724893e-05
R_8_62 n377 PAR_3_0_VDD075NNE 2542.16472581
L_9_62 PAR_1_1_VDD075NNE n378 0.166442382011
R_9_62 n378 PAR_3_0_VDD075NNE 3310.89453983
G0_63 PAR_1_1_VDD075NNE PAR_0_1_VSS PAR_1_1_VDD075NNE PAR_0_1_VSS -0.773059227694
C0_63 PAR_1_1_VDD075NNE PAR_0_1_VSS 2.79556509872e-10
R_1_63 PAR_1_1_VDD075NNE n379 0.0233169272019
C_1_63 n379 PAR_0_1_VSS 1.03797978938e-09
R_2_63 PAR_1_1_VDD075NNE n380 0.012230367046
C_2_63 n380 PAR_0_1_VSS 3.29243114807e-09
L_3_63 PAR_1_1_VDD075NNE n381 2.40371150303e-10
R_3_63 n381 PAR_0_1_VSS 1.70416249893
L_4_63 PAR_1_1_VDD075NNE n382 4.87735949313e-09
R_4_63 n382 PAR_0_1_VSS 5.96142151165
L_5_63 PAR_1_1_VDD075NNE n383 1.79444861324e-07
R_5_63 n383 PAR_0_1_VSS 54.0087923957
R0_64 PAR_1_1_VDD075NNE PAR_0_1_VDD075NNE 0.00251333652937
C0_64 PAR_1_1_VDD075NNE PAR_0_1_VDD075NNE 1.35291655887e-10
L_1_64 PAR_1_1_VDD075NNE n384 2.49735962007e-13
R_1_64 n384 PAR_0_1_VDD075NNE 0.0141624469085
L_2_64 PAR_1_1_VDD075NNE n385 2.24688899483e-13
R_2_64 n385 PAR_0_1_VDD075NNE 0.00602993523829
L_3_64 PAR_1_1_VDD075NNE n386 4.86169227347e-11
R_3_64 n386 PAR_0_1_VDD075NNE 0.652485828915
L_4_64 PAR_1_1_VDD075NNE n387 3.63222692149e-08
R_4_64 n387 PAR_0_1_VDD075NNE 69.0471604938
L_5_64 PAR_1_1_VDD075NNE n388 3.4082475689e-07
R_5_64 n388 PAR_0_1_VDD075NNE 190.334176016
L_6_64 PAR_1_1_VDD075NNE n389 0.00430354581469
R_6_64 n389 PAR_0_1_VDD075NNE 1686.93330388
G0_65 PAR_1_1_VDD075NNE PAR_1_1_VSS PAR_1_1_VDD075NNE PAR_1_1_VSS -0.253644703238
C0_65 PAR_1_1_VDD075NNE PAR_1_1_VSS 1.262840947e-09
R_1_65 PAR_1_1_VDD075NNE n390 0.000391835068868
C_1_65 n390 PAR_1_1_VSS 3.56984280808e-08
R_2_65 PAR_1_1_VDD075NNE n391 0.000261361353173
C_2_65 n391 PAR_1_1_VSS 1.27973557616e-07
R_3_65 PAR_1_1_VDD075NNE n392 0.0094225756093
C_3_65 n392 PAR_1_1_VSS 6.04740244754e-09
R_4_65 PAR_1_1_VDD075NNE n393 0.300021275458
C_4_65 n393 PAR_1_1_VSS 5.0491986807e-10
L_5_65 PAR_1_1_VDD075NNE n394 3.40823165383e-09
R_5_65 n394 PAR_1_1_VSS 4.44201771947
L_6_65 PAR_1_1_VDD075NNE n395 1.03767267262e-07
R_6_65 n395 PAR_1_1_VSS 35.0609171225
G0_66 PAR_1_1_VDD075NNE PAR_0_0_VSS PAR_1_1_VDD075NNE PAR_0_0_VSS -0.244813891346
C0_66 PAR_1_1_VDD075NNE PAR_0_0_VSS 1.95778555909e-10
R_1_66 PAR_1_1_VDD075NNE n396 0.110513187529
C_1_66 n396 PAR_0_0_VSS 1.29638261799e-10
R_2_66 PAR_1_1_VDD075NNE n397 0.25998758292
C_2_66 n397 PAR_0_0_VSS 1.39438463531e-10
L_3_66 PAR_1_1_VDD075NNE n398 7.19394026323e-10
R_3_66 n398 PAR_0_0_VSS 4.70324338878
R_4_66 PAR_1_1_VDD075NNE n399 8.58975341046
C_4_66 n399 PAR_0_0_VSS 4.86917016882e-11
R_5_66 PAR_1_1_VDD075NNE n400 10.3128574594
C_5_66 n400 PAR_0_0_VSS 2.05432037153e-10
L_6_66 PAR_1_1_VDD075NNE n401 2.95920366121e-07
R_6_66 n401 PAR_0_0_VSS 31.0610502445
G0_67 PAR_2_1_VSS PAR_0_0_VDD075NNE PAR_2_1_VSS PAR_0_0_VDD075NNE -1.10040880983
C0_67 PAR_2_1_VSS PAR_0_0_VDD075NNE 2.12740920104e-10
R_1_67 PAR_2_1_VSS n402 0.112967961059
C_1_67 n402 PAR_0_0_VDD075NNE 1.43663510867e-10
L_2_67 PAR_2_1_VSS n403 1.22911830955e-10
R_2_67 n403 PAR_0_0_VDD075NNE 1.72580666328
R_3_67 PAR_2_1_VSS n404 1.55320945232
C_3_67 n404 PAR_0_0_VDD075NNE 8.88675988726e-11
L_4_67 PAR_2_1_VSS n405 1.09101045347e-09
R_4_67 n405 PAR_0_0_VDD075NNE 2.45916935473
L_5_67 PAR_2_1_VSS n406 1.1684052377e-08
R_5_67 n406 PAR_0_0_VDD075NNE 9.21070325868
L_6_67 PAR_2_1_VSS n407 1.23277141284e-06
R_6_67 n407 PAR_0_0_VDD075NNE 173.643772785
R0_68 PAR_2_1_VSS PAR_1_0_VSS 0.152687431263
C0_68 PAR_2_1_VSS PAR_1_0_VSS 2.29364456716e-10
R_1_68 PAR_2_1_VSS n408 0.368500385053
C_1_68 n408 PAR_1_0_VSS 9.59077410721e-11
R_2_68 PAR_2_1_VSS n409 0.616884228119
C_2_68 n409 PAR_1_0_VSS 2.29510880391e-10
R_3_68 PAR_2_1_VSS n410 0.172965703228
C_3_68 n410 PAR_1_0_VSS 2.01669609331e-09
R_4_68 PAR_2_1_VSS n411 1.18975131117
C_4_68 n411 PAR_1_0_VSS 7.3321038047e-10
R_5_68 PAR_2_1_VSS n412 0.822579974094
C_5_68 n412 PAR_1_0_VSS 2.3471623555e-09
L_6_68 PAR_2_1_VSS n413 2.9508647975e-08
R_6_68 n413 PAR_1_0_VSS 3.11116804767
G0_69 PAR_2_1_VSS PAR_1_0_VDD075NNE PAR_2_1_VSS PAR_1_0_VDD075NNE -0.448121487887
C0_69 PAR_2_1_VSS PAR_1_0_VDD075NNE 1.90885012332e-10
R_1_69 PAR_2_1_VSS n414 0.156291171252
C_1_69 n414 PAR_1_0_VDD075NNE 1.15048890322e-10
R_2_69 PAR_2_1_VSS n415 1.96616548562
C_2_69 n415 PAR_1_0_VDD075NNE 8.28155254005e-11
L_3_69 PAR_2_1_VSS n416 1.29439824609e-09
R_3_69 n416 PAR_1_0_VDD075NNE 2.98064492181
L_4_69 PAR_2_1_VSS n417 1.13161574972e-08
R_4_69 n417 PAR_1_0_VDD075NNE 9.34516014731
L_5_69 PAR_2_1_VSS n418 1.21849983825e-06
R_5_69 n418 PAR_1_0_VDD075NNE 178.05106625
R0_70 PAR_2_1_VSS PAR_2_0_VSS 0.0106959429064
C0_70 PAR_2_1_VSS PAR_2_0_VSS 1.6116549934e-10
L_1_70 PAR_2_1_VSS n419 3.81363550737e-13
R_1_70 n419 PAR_2_0_VSS 0.0171332931072
L_2_70 PAR_2_1_VSS n420 3.74395825776e-12
R_2_70 n420 PAR_2_0_VSS 0.0757375512977
R_3_70 PAR_2_1_VSS n421 0.242698427735
C_3_70 n421 PAR_2_0_VSS 1.65314068356e-09
R_4_70 PAR_2_1_VSS n422 1.10805119581
C_4_70 n422 PAR_2_0_VSS 1.36178042759e-09
L_5_70 PAR_2_1_VSS n423 6.55959708566e-08
R_5_70 n423 PAR_2_0_VSS 6.43573494746
G0_71 PAR_2_1_VSS PAR_2_0_VDD075NNE PAR_2_1_VSS PAR_2_0_VDD075NNE -0.442083542575
C0_71 PAR_2_1_VSS PAR_2_0_VDD075NNE 1.90374770477e-10
R_1_71 PAR_2_1_VSS n424 0.0346321120952
C_1_71 n424 PAR_2_0_VDD075NNE 6.49418052238e-10
R_2_71 PAR_2_1_VSS n425 0.11304264254
C_2_71 n425 PAR_2_0_VDD075NNE 3.96579774591e-10
R_3_71 PAR_2_1_VSS n426 1.5507238106
C_3_71 n426 PAR_2_0_VDD075NNE 9.80392623357e-11
L_4_71 PAR_2_1_VSS n427 1.38916572e-09
R_4_71 n427 PAR_2_0_VDD075NNE 2.99232881891
L_5_71 PAR_2_1_VSS n428 1.23753467909e-08
R_5_71 n428 PAR_2_0_VDD075NNE 9.74558393684
L_6_71 PAR_2_1_VSS n429 1.41626073577e-06
R_6_71 n429 PAR_2_0_VDD075NNE 189.211327843
R0_72 PAR_2_1_VSS PAR_3_0_VSS 0.149240573355
C0_72 PAR_2_1_VSS PAR_3_0_VSS 2.36141284545e-10
R_1_72 PAR_2_1_VSS n430 0.0613671510052
C_1_72 n430 PAR_3_0_VSS 7.38014297137e-10
R_2_72 PAR_2_1_VSS n431 0.0964463019228
C_2_72 n431 PAR_3_0_VSS 1.46630411914e-09
R_3_72 PAR_2_1_VSS n432 0.0424767636853
C_3_72 n432 PAR_3_0_VSS 6.8619743327e-09
R_4_72 PAR_2_1_VSS n433 0.136476286997
C_4_72 n433 PAR_3_0_VSS 4.46464458877e-09
R_5_72 PAR_2_1_VSS n434 0.316586204092
C_5_72 n434 PAR_3_0_VSS 3.77743840474e-09
R_6_72 PAR_2_1_VSS n435 1.7562133656
C_6_72 n435 PAR_3_0_VSS 5.60167231959e-09
G0_73 PAR_2_1_VSS PAR_3_0_VDD075NNE PAR_2_1_VSS PAR_3_0_VDD075NNE -1.46159685663
C0_73 PAR_2_1_VSS PAR_3_0_VDD075NNE 2.5113252457e-10
R_1_73 PAR_2_1_VSS n436 0.0498952068321
C_1_73 n436 PAR_3_0_VDD075NNE 3.76748513078e-10
R_2_73 PAR_2_1_VSS n437 0.36496420488
C_2_73 n437 PAR_3_0_VDD075NNE 1.16107842922e-10
R_3_73 PAR_2_1_VSS n438 0.748715065681
C_3_73 n438 PAR_3_0_VDD075NNE 2.34458048631e-10
L_4_73 PAR_2_1_VSS n439 3.68661881293e-10
R_4_73 n439 PAR_3_0_VDD075NNE 0.832766427016
L_5_73 PAR_2_1_VSS n440 4.78386621445e-09
R_5_73 n440 PAR_3_0_VDD075NNE 4.00909583461
L_6_73 PAR_2_1_VSS n441 4.86673611365e-07
R_6_73 n441 PAR_3_0_VDD075NNE 88.1277872207
G0_74 PAR_2_1_VSS PAR_0_1_VSS PAR_2_1_VSS PAR_0_1_VSS -9.80413987748
C0_74 PAR_2_1_VSS PAR_0_1_VSS 2.71446111869e-10
R_1_74 PAR_2_1_VSS n442 0.0923304983259
C_1_74 n442 PAR_0_1_VSS 3.63135785965e-10
R_2_74 PAR_2_1_VSS n443 0.0403498679463
C_2_74 n443 PAR_0_1_VSS 5.86997570019e-09
L_3_74 PAR_2_1_VSS n444 5.22172706626e-11
R_3_74 n444 PAR_0_1_VSS 0.125476320075
L_4_74 PAR_2_1_VSS n445 6.48095938752e-10
R_4_74 n445 PAR_0_1_VSS 0.556548302949
L_5_74 PAR_2_1_VSS n446 7.95981952e-08
R_5_74 n446 PAR_0_1_VSS 11.8849434451
G0_75 PAR_2_1_VSS PAR_0_1_VDD075NNE PAR_2_1_VSS PAR_0_1_VDD075NNE -1.00606523493
C0_75 PAR_2_1_VSS PAR_0_1_VDD075NNE 2.54335041004e-10
R_1_75 PAR_2_1_VSS n447 0.0559834082259
C_1_75 n447 PAR_0_1_VDD075NNE 2.12658627115e-10
R_2_75 PAR_2_1_VSS n448 1.85239512647
C_2_75 n448 PAR_0_1_VDD075NNE 9.22984321103e-11
L_3_75 PAR_2_1_VSS n449 3.6760382491e-10
R_3_75 n449 PAR_0_1_VDD075NNE 1.28092396734
L_4_75 PAR_2_1_VSS n450 4.53902527545e-09
R_4_75 n450 PAR_0_1_VDD075NNE 4.75371025137
L_5_75 PAR_2_1_VSS n451 3.12815929229e-07
R_5_75 n451 PAR_0_1_VDD075NNE 66.5921913862
R0_76 PAR_2_1_VSS PAR_1_1_VSS 0.00236819086842
C0_76 PAR_2_1_VSS PAR_1_1_VSS 7.3812807653e-12
L_1_76 PAR_2_1_VSS n452 1.62404597436e-13
R_1_76 n452 PAR_1_1_VSS 0.00512028666468
L_2_76 PAR_2_1_VSS n453 1.81327095893e-11
R_2_76 n453 PAR_1_1_VSS 0.213515297929
R_3_76 PAR_2_1_VSS n454 0.146565118376
C_3_76 n454 PAR_1_1_VSS 1.17552151091e-09
L_4_76 PAR_2_1_VSS n455 5.64743354412e-11
R_4_76 n455 PAR_1_1_VSS 0.118500853797
L_5_76 PAR_2_1_VSS n456 7.42241793115e-10
R_5_76 n456 PAR_1_1_VSS 0.568321275821
L_6_76 PAR_2_1_VSS n457 9.87662108924e-08
R_6_76 n457 PAR_1_1_VSS 12.3776596658
G0_77 PAR_2_1_VSS PAR_1_1_VDD075NNE PAR_2_1_VSS PAR_1_1_VDD075NNE -0.420604356511
C0_77 PAR_2_1_VSS PAR_1_1_VDD075NNE 2.27250566232e-10
R_1_77 PAR_2_1_VSS n458 0.0231509476069
C_1_77 n458 PAR_1_1_VDD075NNE 6.92036749781e-10
R_2_77 PAR_2_1_VSS n459 0.0108738266183
C_2_77 n459 PAR_1_1_VDD075NNE 3.37576823952e-09
R_3_77 PAR_2_1_VSS n460 1.50250693842
C_3_77 n460 PAR_1_1_VDD075NNE 9.57251327333e-11
L_4_77 PAR_2_1_VSS n461 1.55881078544e-09
R_4_77 n461 PAR_1_1_VDD075NNE 3.37550552478
L_5_77 PAR_2_1_VSS n462 1.06198230346e-08
R_5_77 n462 PAR_1_1_VDD075NNE 8.48324341556
L_6_77 PAR_2_1_VSS n463 1.15120161789e-06
R_6_77 n463 PAR_1_1_VDD075NNE 154.487989911
G0_78 PAR_2_1_VSS PAR_0_0_VSS PAR_2_1_VSS PAR_0_0_VSS -0.444473380376
C0_78 PAR_2_1_VSS PAR_0_0_VSS 2.06681851529e-10
R_1_78 PAR_2_1_VSS n464 0.129827177889
C_1_78 n464 PAR_0_0_VSS 2.93460323283e-10
R_2_78 PAR_2_1_VSS n465 0.631378128919
C_2_78 n465 PAR_0_0_VSS 1.98406939103e-10
R_3_78 PAR_2_1_VSS n466 0.134252698215
C_3_78 n466 PAR_0_0_VSS 2.08062080931e-09
R_4_78 PAR_2_1_VSS n467 0.245813474304
C_4_78 n467 PAR_0_0_VSS 1.74315825269e-09
R_5_78 PAR_2_1_VSS n468 0.677550716087
C_5_78 n468 PAR_0_0_VSS 3.14095688067e-09
L_6_78 PAR_2_1_VSS n469 2.13896929843e-08
R_6_78 n469 PAR_0_0_VSS 2.24982361541
G0_79 PAR_2_1_VDD075NNE PAR_0_0_VDD075NNE PAR_2_1_VDD075NNE PAR_0_0_VDD075NNE -7.54820025444
C0_79 PAR_2_1_VDD075NNE PAR_0_0_VDD075NNE 1.30962909421e-10
R_1_79 PAR_2_1_VDD075NNE n470 0.180320472727
C_1_79 n470 PAR_0_0_VDD075NNE 1.31301410581e-10
L_2_79 PAR_2_1_VDD075NNE n471 7.85537945514e-12
R_2_79 n471 PAR_0_0_VDD075NNE 0.150319814345
R_3_79 PAR_2_1_VDD075NNE n472 0.596372729344
C_3_79 n472 PAR_0_0_VDD075NNE 2.16605872899e-10
L_4_79 PAR_2_1_VDD075NNE n473 3.92587830823e-10
R_4_79 n473 PAR_0_0_VDD075NNE 1.30882474319
R_5_79 PAR_2_1_VDD075NNE n474 3.07231748274
C_5_79 n474 PAR_0_0_VDD075NNE 2.70090167039e-10
L_6_79 PAR_2_1_VDD075NNE n475 1.53976088641e-08
R_6_79 n475 PAR_0_0_VDD075NNE 7.56494985355
R_7_79 PAR_2_1_VDD075NNE n476 4398.36978277
C_7_79 n476 PAR_0_0_VDD075NNE 2.53302116814e-10
G0_80 PAR_2_1_VDD075NNE PAR_1_0_VSS PAR_2_1_VDD075NNE PAR_1_0_VSS -0.129938043888
C0_80 PAR_2_1_VDD075NNE PAR_1_0_VSS 2.28073258242e-10
R_1_80 PAR_2_1_VDD075NNE n477 0.0791856417884
C_1_80 n477 PAR_1_0_VSS 2.06539933101e-10
R_2_80 PAR_2_1_VDD075NNE n478 0.316530459863
C_2_80 n478 PAR_1_0_VSS 1.2741576863e-10
L_3_80 PAR_2_1_VDD075NNE n479 1.26042881362e-09
R_3_80 n479 PAR_1_0_VSS 9.42694382908
R_4_80 PAR_2_1_VDD075NNE n480 11.1205396224
C_4_80 n480 PAR_1_0_VSS 4.26718520982e-11
R_5_80 PAR_2_1_VDD075NNE n481 9.73209559448
C_5_80 n481 PAR_1_0_VSS 1.7937339892e-10
L_6_80 PAR_2_1_VDD075NNE n482 4.10741540531e-07
R_6_80 n482 PAR_1_0_VSS 41.9126752929
G0_81 PAR_2_1_VDD075NNE PAR_1_0_VDD075NNE PAR_2_1_VDD075NNE PAR_1_0_VDD075NNE -0.21668786075
C0_81 PAR_2_1_VDD075NNE PAR_1_0_VDD075NNE 1.53439360025e-10
L_1_81 PAR_2_1_VDD075NNE n483 4.34372204984e-12
R_1_81 n483 PAR_1_0_VDD075NNE 0.196354697956
L_2_81 PAR_2_1_VDD075NNE n484 1.88855695206e-11
R_2_81 n484 PAR_1_0_VDD075NNE 0.35463874283
R_3_81 PAR_2_1_VDD075NNE n485 5.04256787985
C_3_81 n485 PAR_1_0_VDD075NNE 3.31921885934e-11
L_4_81 PAR_2_1_VDD075NNE n486 7.40301183002e-09
R_4_81 n486 PAR_1_0_VDD075NNE 10.6831760769
R_5_81 PAR_2_1_VDD075NNE n487 54.4182085806
C_5_81 n487 PAR_1_0_VDD075NNE 4.26710845559e-11
G0_82 PAR_2_1_VDD075NNE PAR_2_0_VSS PAR_2_1_VDD075NNE PAR_2_0_VSS -0.0126964466272
C0_82 PAR_2_1_VDD075NNE PAR_2_0_VSS 2.47510994211e-10
R_1_82 PAR_2_1_VDD075NNE n488 0.00686488524998
C_1_82 n488 PAR_2_0_VSS 2.41694347154e-09
R_2_82 PAR_2_1_VDD075NNE n489 0.0197062661739
C_2_82 n489 PAR_2_0_VSS 1.94340140455e-09
R_3_82 PAR_2_1_VDD075NNE n490 0.791170576539
C_3_82 n490 PAR_2_0_VSS 9.85957460008e-11
R_4_82 PAR_2_1_VDD075NNE n491 10.0295202363
C_4_82 n491 PAR_2_0_VSS 4.18772979616e-11
R_5_82 PAR_2_1_VDD075NNE n492 17.3624164263
C_5_82 n492 PAR_2_0_VSS 9.023777555e-11
L_6_82 PAR_2_1_VDD075NNE n493 7.77037255e-07
R_6_82 n493 PAR_2_0_VSS 78.7621678282
R0_83 PAR_2_1_VDD075NNE PAR_2_0_VDD075NNE 0.00812339780322
C0_83 PAR_2_1_VDD075NNE PAR_2_0_VDD075NNE 1.69660630776e-10
L_1_83 PAR_2_1_VDD075NNE n494 2.59310925316e-13
R_1_83 n494 PAR_2_0_VDD075NNE 0.0128133338167
L_2_83 PAR_2_1_VDD075NNE n495 1.78039344811e-12
R_2_83 n495 PAR_2_0_VDD075NNE 0.0429147580647
L_3_83 PAR_2_1_VDD075NNE n496 4.21230264586e-10
R_3_83 n496 PAR_2_0_VDD075NNE 3.83261548904
L_4_83 PAR_2_1_VDD075NNE n497 3.04291638363e-08
R_4_83 n497 PAR_2_0_VDD075NNE 64.6677705308
L_5_83 PAR_2_1_VDD075NNE n498 3.24654769142e-07
R_5_83 n498 PAR_2_0_VDD075NNE 194.304756828
L_6_83 PAR_2_1_VDD075NNE n499 0.00655716940797
R_6_83 n499 PAR_2_0_VDD075NNE 1017.99037014
G0_84 PAR_2_1_VDD075NNE PAR_3_0_VSS PAR_2_1_VDD075NNE PAR_3_0_VSS -0.830216554798
C0_84 PAR_2_1_VDD075NNE PAR_3_0_VSS 2.83696689407e-10
R_1_84 PAR_2_1_VDD075NNE n500 0.021433058846
C_1_84 n500 PAR_3_0_VSS 7.78265535282e-10
R_2_84 PAR_2_1_VDD075NNE n501 0.121154212225
C_2_84 n501 PAR_3_0_VSS 3.73938188837e-10
L_3_84 PAR_2_1_VDD075NNE n502 1.91124627309e-10
R_3_84 n502 PAR_3_0_VSS 1.20450500121
R_4_84 PAR_2_1_VDD075NNE n503 3.20307417523
C_4_84 n503 PAR_3_0_VSS 1.80333301328e-10
R_5_84 PAR_2_1_VDD075NNE n504 4.4810947884
C_5_84 n504 PAR_3_0_VSS 2.57336407093e-10
R_6_84 PAR_2_1_VDD075NNE n505 22.4171763095
C_6_84 n505 PAR_3_0_VSS 4.37159105099e-10
G0_85 PAR_2_1_VDD075NNE PAR_3_0_VDD075NNE PAR_2_1_VDD075NNE PAR_3_0_VDD075NNE -4.15013168549
C0_85 PAR_2_1_VDD075NNE PAR_3_0_VDD075NNE 1.93438967944e-10
R_1_85 PAR_2_1_VDD075NNE n506 0.0225266027859
C_1_85 n506 PAR_3_0_VDD075NNE 1.78490019315e-10
L_2_85 PAR_2_1_VDD075NNE n507 3.133848976e-12
R_2_85 n507 PAR_3_0_VDD075NNE 0.106571076604
L_3_85 PAR_2_1_VDD075NNE n508 2.56865392985e-11
R_3_85 n508 PAR_3_0_VDD075NNE 0.425576377756
L_4_85 PAR_2_1_VDD075NNE n509 1.05589913249e-09
R_4_85 n509 PAR_3_0_VDD075NNE 7.48927847255
L_5_85 PAR_2_1_VDD075NNE n510 6.66756329546e-09
R_5_85 n510 PAR_3_0_VDD075NNE 21.8321699064
L_6_85 PAR_2_1_VDD075NNE n511 3.44448722688e-08
R_6_85 n511 PAR_3_0_VDD075NNE 48.2931514883
L_7_85 PAR_2_1_VDD075NNE n512 1.88443830515e-07
R_7_85 n512 PAR_3_0_VDD075NNE 117.041160573
R_8_85 PAR_2_1_VDD075NNE n513 2646.24034048
C_8_85 n513 PAR_3_0_VDD075NNE 3.04953075588e-12
G0_86 PAR_2_1_VDD075NNE PAR_0_1_VSS PAR_2_1_VDD075NNE PAR_0_1_VSS -0.870711811573
C0_86 PAR_2_1_VDD075NNE PAR_0_1_VSS 2.79287075932e-10
R_1_86 PAR_2_1_VDD075NNE n514 0.110871414915
C_1_86 n514 PAR_0_1_VSS 1.30454270857e-10
R_2_86 PAR_2_1_VDD075NNE n515 3.6839852843
C_2_86 n515 PAR_0_1_VSS 2.97418530543e-11
L_3_86 PAR_2_1_VDD075NNE n516 3.81283294949e-10
R_3_86 n516 PAR_0_1_VSS 1.42723614346
L_4_86 PAR_2_1_VDD075NNE n517 5.92090505931e-09
R_4_86 n517 PAR_0_1_VSS 6.34478155652
L_5_86 PAR_2_1_VDD075NNE n518 3.57175187716e-07
R_5_86 n518 PAR_0_1_VSS 80.3401565809
G0_87 PAR_2_1_VDD075NNE PAR_0_1_VDD075NNE PAR_2_1_VDD075NNE PAR_0_1_VDD075NNE -8.9525910855
C0_87 PAR_2_1_VDD075NNE PAR_0_1_VDD075NNE 1.6496656615e-10
R_1_87 PAR_2_1_VDD075NNE n519 0.16113164588
C_1_87 n519 PAR_0_1_VDD075NNE 1.55040880794e-10
L_2_87 PAR_2_1_VDD075NNE n520 7.41021725101e-12
R_2_87 n520 PAR_0_1_VDD075NNE 0.120636506323
R_3_87 PAR_2_1_VDD075NNE n521 0.414121106974
C_3_87 n521 PAR_0_1_VDD075NNE 2.86107841053e-10
L_4_87 PAR_2_1_VDD075NNE n522 9.34465845127e-10
R_4_87 n522 PAR_0_1_VDD075NNE 1.74515883157
R_5_87 PAR_2_1_VDD075NNE n523 3.01447253439
C_5_87 n523 PAR_0_1_VDD075NNE 4.10981051328e-10
L_6_87 PAR_2_1_VDD075NNE n524 6.36487067626e-08
R_6_87 n524 PAR_0_1_VDD075NNE 11.1862110491
G0_88 PAR_2_1_VDD075NNE PAR_1_1_VSS PAR_2_1_VDD075NNE PAR_1_1_VSS -0.505679854006
C0_88 PAR_2_1_VDD075NNE PAR_1_1_VSS 3.12480547148e-10
R_1_88 PAR_2_1_VDD075NNE n525 0.00533522130307
C_1_88 n525 PAR_1_1_VSS 2.71288316974e-09
R_2_88 PAR_2_1_VDD075NNE n526 0.00401122361203
C_2_88 n526 PAR_1_1_VSS 8.65502519236e-09
R_3_88 PAR_2_1_VDD075NNE n527 0.31397639071
C_3_88 n527 PAR_1_1_VSS 2.36468468581e-10
L_4_88 PAR_2_1_VDD075NNE n528 1.10211761781e-09
R_4_88 n528 PAR_1_1_VSS 2.88790177993
L_5_88 PAR_2_1_VDD075NNE n529 7.47406612476e-09
R_5_88 n529 PAR_1_1_VSS 6.64324271781
L_6_88 PAR_2_1_VDD075NNE n530 7.11692841889e-07
R_6_88 n530 PAR_1_1_VSS 112.627864295
R0_89 PAR_2_1_VDD075NNE PAR_1_1_VDD075NNE 0.0027319737967
C0_89 PAR_2_1_VDD075NNE PAR_1_1_VDD075NNE 1.04907273725e-10
L_1_89 PAR_2_1_VDD075NNE n531 1.41807642042e-13
R_1_89 n531 PAR_1_1_VDD075NNE 0.00851476642069
L_2_89 PAR_2_1_VDD075NNE n532 2.54847786103e-13
R_2_89 n532 PAR_1_1_VDD075NNE 0.0069712953694
L_3_89 PAR_2_1_VDD075NNE n533 1.73111864339e-10
R_3_89 n533 PAR_1_1_VDD075NNE 1.81809878596
L_4_89 PAR_2_1_VDD075NNE n534 2.57590785464e-08
R_4_89 n534 PAR_1_1_VDD075NNE 60.9700382156
L_5_89 PAR_2_1_VDD075NNE n535 2.45619761591e-07
R_5_89 n535 PAR_1_1_VDD075NNE 154.598073113
L_6_89 PAR_2_1_VDD075NNE n536 0.00493158645533
R_6_89 n536 PAR_1_1_VDD075NNE 927.881705499
G0_90 PAR_2_1_VDD075NNE PAR_2_1_VSS PAR_2_1_VDD075NNE PAR_2_1_VSS -0.236711296113
C0_90 PAR_2_1_VDD075NNE PAR_2_1_VSS 9.09410466304e-10
R_1_90 PAR_2_1_VDD075NNE n537 0.000436816359992
C_1_90 n537 PAR_2_1_VSS 3.00497757291e-08
R_2_90 PAR_2_1_VDD075NNE n538 0.000254904368398
C_2_90 n538 PAR_2_1_VSS 1.27793322595e-07
R_3_90 PAR_2_1_VDD075NNE n539 0.00418971260434
C_3_90 n539 PAR_2_1_VSS 1.21511827471e-08
R_4_90 PAR_2_1_VDD075NNE n540 0.409896106533
C_4_90 n540 PAR_2_1_VSS 4.82466528957e-10
L_5_90 PAR_2_1_VDD075NNE n541 4.10523111995e-09
R_5_90 n541 PAR_2_1_VSS 4.58248809972
L_6_90 PAR_2_1_VDD075NNE n542 2.16672799669e-07
R_6_90 n542 PAR_2_1_VSS 54.0855156832
G0_91 PAR_2_1_VDD075NNE PAR_0_0_VSS PAR_2_1_VDD075NNE PAR_0_0_VSS -0.0221966305129
C0_91 PAR_2_1_VDD075NNE PAR_0_0_VSS 2.09582487339e-10
R_1_91 PAR_2_1_VDD075NNE n543 0.120688697792
C_1_91 n543 PAR_0_0_VSS 1.43579729168e-10
R_2_91 PAR_2_1_VDD075NNE n544 7.29301605428
C_2_91 n544 PAR_0_0_VSS 2.08252077072e-10
L_3_91 PAR_2_1_VDD075NNE n545 1.27276740523e-06
R_3_91 n545 PAR_0_0_VSS 45.0518747916
G0_92 PAR_3_1_VSS PAR_0_0_VDD075NNE PAR_3_1_VSS PAR_0_0_VDD075NNE -0.789116954253
C0_92 PAR_3_1_VSS PAR_0_0_VDD075NNE 3.20437384634e-10
R_1_92 PAR_3_1_VSS n546 0.0266624582036
C_1_92 n546 PAR_0_0_VDD075NNE 8.13099251338e-10
L_2_92 PAR_3_1_VSS n547 1.78351956714e-10
R_2_92 n547 PAR_0_0_VDD075NNE 1.33494570402
L_3_92 PAR_3_1_VSS n548 8.90763515634e-08
R_3_92 n548 PAR_0_0_VDD075NNE 24.9857446546
R0_93 PAR_3_1_VSS PAR_1_0_VSS 10.1794038071
C0_93 PAR_3_1_VSS PAR_1_0_VSS 3.00552009455e-10
R_1_93 PAR_3_1_VSS n549 0.0531057031121
C_1_93 n549 PAR_1_0_VSS 5.46503135897e-10
R_2_93 PAR_3_1_VSS n550 0.0824323746149
C_2_93 n550 PAR_1_0_VSS 1.20476500053e-09
R_3_93 PAR_3_1_VSS n551 0.279025022282
C_3_93 n551 PAR_1_0_VSS 8.51680557461e-10
R_4_93 PAR_3_1_VSS n552 0.16881652273
C_4_93 n552 PAR_1_0_VSS 3.32689362343e-09
R_5_93 PAR_3_1_VSS n553 0.119233074555
C_5_93 n553 PAR_1_0_VSS 2.11865131361e-08
R_6_93 PAR_3_1_VSS n554 0.222642303722
C_6_93 n554 PAR_1_0_VSS 3.82230537087e-08
G0_94 PAR_3_1_VSS PAR_1_0_VDD075NNE PAR_3_1_VSS PAR_1_0_VDD075NNE -0.524867141847
C0_94 PAR_3_1_VSS PAR_1_0_VDD075NNE 2.31677825034e-10
R_1_94 PAR_3_1_VSS n555 0.0301823518949
C_1_94 n555 PAR_1_0_VDD075NNE 4.57571143101e-10
R_2_94 PAR_3_1_VSS n556 0.147955080033
C_2_94 n556 PAR_1_0_VDD075NNE 2.40876950931e-10
L_3_94 PAR_3_1_VSS n557 2.93606431566e-10
R_3_94 n557 PAR_1_0_VDD075NNE 2.34877315743
R_4_94 PAR_3_1_VSS n558 8.09671306423
C_4_94 n558 PAR_1_0_VDD075NNE 6.29066599421e-11
L_5_94 PAR_3_1_VSS n559 2.3310742748e-08
R_5_94 n559 PAR_1_0_VDD075NNE 10.089497697
R_6_94 PAR_3_1_VSS n560 29.7340751384
C_6_94 n560 PAR_1_0_VDD075NNE 2.93218898527e-10
R0_95 PAR_3_1_VSS PAR_2_0_VSS 0.144942557526
C0_95 PAR_3_1_VSS PAR_2_0_VSS 2.80698182873e-10
R_1_95 PAR_3_1_VSS n561 0.0659427133884
C_1_95 n561 PAR_2_0_VSS 2.84137556002e-10
R_2_95 PAR_3_1_VSS n562 0.295008755659
C_2_95 n562 PAR_2_0_VSS 4.01371255993e-10
R_3_95 PAR_3_1_VSS n563 0.268131098821
C_3_95 n563 PAR_2_0_VSS 1.77382309753e-09
R_4_95 PAR_3_1_VSS n564 0.506465976256
C_4_95 n564 PAR_2_0_VSS 1.67594448141e-09
R_5_95 PAR_3_1_VSS n565 0.203893369306
C_5_95 n565 PAR_2_0_VSS 1.19842308223e-08
R_6_95 PAR_3_1_VSS n566 0.384460721065
C_6_95 n566 PAR_2_0_VSS 2.2565627315e-08
G0_96 PAR_3_1_VSS PAR_2_0_VDD075NNE PAR_3_1_VSS PAR_2_0_VDD075NNE -0.030256187636
C0_96 PAR_3_1_VSS PAR_2_0_VDD075NNE 3.61240256384e-10
R_1_96 PAR_3_1_VSS n567 0.0414455031945
C_1_96 n567 PAR_2_0_VDD075NNE 6.41748545259e-10
R_2_96 PAR_3_1_VSS n568 11.7720385958
C_2_96 n568 PAR_2_0_VDD075NNE 4.30015365872e-11
L_3_96 PAR_3_1_VSS n569 1.46379998115e-07
R_3_96 n569 PAR_2_0_VDD075NNE 33.0510853596
R0_97 PAR_3_1_VSS PAR_3_0_VSS 0.0113160692565
C0_97 PAR_3_1_VSS PAR_3_0_VSS 2.77872348417e-10
L_1_97 PAR_3_1_VSS n570 1.22775168185e-13
R_1_97 n570 PAR_3_0_VSS 0.00774428647797
R_2_97 PAR_3_1_VSS n571 0.0145181990741
C_2_97 n571 PAR_3_0_VSS 7.2820762235e-09
R_3_97 PAR_3_1_VSS n572 0.0456007668458
C_3_97 n572 PAR_3_0_VSS 5.75706561358e-09
R_4_97 PAR_3_1_VSS n573 0.0555975346138
C_4_97 n573 PAR_3_0_VSS 1.30572498067e-08
R_5_97 PAR_3_1_VSS n574 0.0558394664783
C_5_97 n574 PAR_3_0_VSS 3.11565805362e-08
R_6_97 PAR_3_1_VSS n575 0.196028712731
C_6_97 n575 PAR_3_0_VSS 5.67715829254e-08
G0_98 PAR_3_1_VSS PAR_3_0_VDD075NNE PAR_3_1_VSS PAR_3_0_VDD075NNE -0.603407304343
C0_98 PAR_3_1_VSS PAR_3_0_VDD075NNE 4.46827357085e-10
R_1_98 PAR_3_1_VSS n576 0.0109100182297
C_1_98 n576 PAR_3_0_VDD075NNE 2.88874346388e-09
L_2_98 PAR_3_1_VSS n577 8.17076808638e-09
R_2_98 n577 PAR_3_0_VDD075NNE 19.0974268729
L_3_98 PAR_3_1_VSS n578 1.96670233836e-09
R_3_98 n578 PAR_3_0_VDD075NNE 1.81473634629
R0_99 PAR_3_1_VSS PAR_0_1_VSS 4320.69850391
C0_99 PAR_3_1_VSS PAR_0_1_VSS 4.42286958251e-10
R_1_99 PAR_3_1_VSS n579 0.0314582065141
C_1_99 n579 PAR_0_1_VSS 2.08010114462e-09
R_2_99 PAR_3_1_VSS n580 0.0242379745075
C_2_99 n580 PAR_0_1_VSS 8.98051581253e-09
R_3_99 PAR_3_1_VSS n581 3.42630193568
C_3_99 n581 PAR_0_1_VSS 8.11543231097e-10
G0_100 PAR_3_1_VSS PAR_0_1_VDD075NNE PAR_3_1_VSS PAR_0_1_VDD075NNE -2.09029575091
C0_100 PAR_3_1_VSS PAR_0_1_VDD075NNE 4.69512226132e-10
R_1_100 PAR_3_1_VSS n582 0.0210465734597
C_1_100 n582 PAR_0_1_VDD075NNE 1.10036190532e-09
L_2_100 PAR_3_1_VSS n583 7.65108355809e-11
R_2_100 n583 PAR_0_1_VDD075NNE 0.479219415229
L_3_100 PAR_3_1_VSS n584 1.30952978366e-05
R_3_100 n584 PAR_0_1_VDD075NNE 280.194471155
R0_101 PAR_3_1_VSS PAR_1_1_VSS 11.7483408668
C0_101 PAR_3_1_VSS PAR_1_1_VSS 4.85353463226e-10
R_1_101 PAR_3_1_VSS n585 0.0350989824917
C_1_101 n585 PAR_1_1_VSS 2.06229488121e-09
R_2_101 PAR_3_1_VSS n586 0.0189970485357
C_2_101 n586 PAR_1_1_VSS 1.17669157544e-08
R_3_101 PAR_3_1_VSS n587 3.52488210309
C_3_101 n587 PAR_1_1_VSS 1.04187699333e-09
G0_102 PAR_3_1_VSS PAR_1_1_VDD075NNE PAR_3_1_VSS PAR_1_1_VDD075NNE -1.22104628579
C0_102 PAR_3_1_VSS PAR_1_1_VDD075NNE 4.15857609046e-10
R_1_102 PAR_3_1_VSS n588 0.0248382309255
C_1_102 n588 PAR_1_1_VDD075NNE 8.97590116166e-10
L_2_102 PAR_3_1_VSS n589 1.38131303095e-10
R_2_102 n589 PAR_1_1_VDD075NNE 0.821728217054
L_3_102 PAR_3_1_VSS n590 8.61624150011e-06
R_3_102 n590 PAR_1_1_VDD075NNE 243.967235736
R0_103 PAR_3_1_VSS PAR_2_1_VSS 0.00213041546035
C0_103 PAR_3_1_VSS PAR_2_1_VSS 4.8667555647e-11
L_1_103 PAR_3_1_VSS n591 1.93336715515e-13
R_1_103 n591 PAR_2_1_VSS 0.00612930972231
R_2_103 PAR_3_1_VSS n592 0.056782055564
C_2_103 n592 PAR_2_1_VSS 3.61167894149e-09
R_3_103 PAR_3_1_VSS n593 0.0736975560292
C_3_103 n593 PAR_2_1_VSS 5.02613252506e-09
L_4_103 PAR_3_1_VSS n594 1.70401606479e-09
R_4_103 n594 PAR_2_1_VSS 0.614089975705
R_5_103 PAR_3_1_VSS n595 1.22759781566
C_5_103 n595 PAR_2_1_VSS 6.29595057487e-09
C0_104 PAR_3_1_VSS PAR_2_1_VDD075NNE 1.06787354519e-09
R_1_104 PAR_3_1_VSS n596 0.00291343790278
C_1_104 n596 PAR_2_1_VDD075NNE 1.1484773479e-08
R0_105 PAR_3_1_VSS PAR_0_0_VSS 23.3543448958
C0_105 PAR_3_1_VSS PAR_0_0_VSS 2.25633393776e-10
R_1_105 PAR_3_1_VSS n597 0.0583109273694
C_1_105 n597 PAR_0_0_VSS 8.44733762603e-10
R_2_105 PAR_3_1_VSS n598 0.0625429655929
C_2_105 n598 PAR_0_0_VSS 1.847020011e-09
R_3_105 PAR_3_1_VSS n599 0.143469081057
C_3_105 n599 PAR_0_0_VSS 1.7448728889e-09
R_4_105 PAR_3_1_VSS n600 0.0923373051095
C_4_105 n600 PAR_0_0_VSS 6.10227107754e-09
R_5_105 PAR_3_1_VSS n601 0.104756840108
C_5_105 n601 PAR_0_0_VSS 2.64814063198e-08
R_6_105 PAR_3_1_VSS n602 0.172570298334
C_6_105 n602 PAR_0_0_VSS 4.93260987031e-08
G0_106 PAR_3_1_VDD075NNE PAR_0_0_VDD075NNE PAR_3_1_VDD075NNE PAR_0_0_VDD075NNE -8.75313032572
C0_106 PAR_3_1_VDD075NNE PAR_0_0_VDD075NNE 1.5158171148e-10
R_1_106 PAR_3_1_VDD075NNE n603 0.0179202323523
C_1_106 n603 PAR_0_0_VDD075NNE 1.49073710556e-10
L_2_106 PAR_3_1_VDD075NNE n604 3.83794756911e-12
R_2_106 n604 PAR_0_0_VDD075NNE 0.136245890747
L_3_106 PAR_3_1_VDD075NNE n605 3.6554902141e-11
R_3_106 n605 PAR_0_0_VDD075NNE 0.737321983667
L_4_106 PAR_3_1_VDD075NNE n606 4.37136433473e-09
R_4_106 n606 PAR_0_0_VDD075NNE 32.6022698861
L_5_106 PAR_3_1_VDD075NNE n607 2.25563020032e-08
R_5_106 n607 PAR_0_0_VDD075NNE 63.9039628285
L_6_106 PAR_3_1_VDD075NNE n608 1.11844467367e-07
R_6_106 n608 PAR_0_0_VDD075NNE 139.175788652
L_7_106 PAR_3_1_VDD075NNE n609 4.63764392438e-07
R_7_106 n609 PAR_0_0_VDD075NNE 284.793875969
G0_107 PAR_3_1_VDD075NNE PAR_1_0_VSS PAR_3_1_VDD075NNE PAR_1_0_VSS -0.945772909985
C0_107 PAR_3_1_VDD075NNE PAR_1_0_VSS 2.0432634531e-10
R_1_107 PAR_3_1_VDD075NNE n610 0.0526760386646
C_1_107 n610 PAR_1_0_VSS 1.43216372276e-10
L_2_107 PAR_3_1_VDD075NNE n611 1.11925484695e-10
R_2_107 n611 PAR_1_0_VSS 1.33477713244
L_3_107 PAR_3_1_VDD075NNE n612 1.02550805009e-09
R_3_107 n612 PAR_1_0_VSS 5.83082036014
R_4_107 PAR_3_1_VDD075NNE n613 8.59886849549
C_4_107 n613 PAR_1_0_VSS 4.10049938513e-11
R_5_107 PAR_3_1_VDD075NNE n614 11.2421008421
C_5_107 n614 PAR_1_0_VSS 1.45168815883e-10
L_6_107 PAR_3_1_VDD075NNE n615 3.81222579823e-07
R_6_107 n615 PAR_1_0_VSS 39.8696771718
G0_108 PAR_3_1_VDD075NNE PAR_1_0_VDD075NNE PAR_3_1_VDD075NNE PAR_1_0_VDD075NNE -8.98505765148
C0_108 PAR_3_1_VDD075NNE PAR_1_0_VDD075NNE 1.29369341128e-10
R_1_108 PAR_3_1_VDD075NNE n616 0.165908486623
C_1_108 n616 PAR_1_0_VDD075NNE 1.71854491337e-10
L_2_108 PAR_3_1_VDD075NNE n617 8.01794675361e-12
R_2_108 n617 PAR_1_0_VDD075NNE 0.138257300617
R_3_108 PAR_3_1_VDD075NNE n618 0.505467211762
C_3_108 n618 PAR_1_0_VDD075NNE 3.16309457935e-10
L_4_108 PAR_3_1_VDD075NNE n619 3.05707446424e-10
R_4_108 n619 PAR_1_0_VDD075NNE 0.77459906086
R_5_108 PAR_3_1_VDD075NNE n620 1.05796268711
C_5_108 n620 PAR_1_0_VDD075NNE 8.79644942854e-10
L_6_108 PAR_3_1_VDD075NNE n621 3.92773565083e-09
R_6_108 n621 PAR_1_0_VDD075NNE 2.16771875173
R_7_108 PAR_3_1_VDD075NNE n622 29.3618249138
C_7_108 n622 PAR_1_0_VDD075NNE 3.12318461428e-10
G0_109 PAR_3_1_VDD075NNE PAR_2_0_VSS PAR_3_1_VDD075NNE PAR_2_0_VSS -0.00203223556673
C0_109 PAR_3_1_VDD075NNE PAR_2_0_VSS 2.30202413921e-10
R_1_109 PAR_3_1_VDD075NNE n623 0.613430890044
C_1_109 n623 PAR_2_0_VSS 4.95613421576e-11
R_2_109 PAR_3_1_VDD075NNE n624 8.85729628809
C_2_109 n624 PAR_2_0_VSS 6.39597320479e-11
L_3_109 PAR_3_1_VDD075NNE n625 8.19570180592e-05
R_3_109 n625 PAR_2_0_VSS 492.06818571
G0_110 PAR_3_1_VDD075NNE PAR_2_0_VDD075NNE PAR_3_1_VDD075NNE PAR_2_0_VDD075NNE -0.528533363668
C0_110 PAR_3_1_VDD075NNE PAR_2_0_VDD075NNE 1.9370819442e-10
L_1_110 PAR_3_1_VDD075NNE n626 5.50952126891e-12
R_1_110 n626 PAR_2_0_VDD075NNE 0.191751227896
L_2_110 PAR_3_1_VDD075NNE n627 2.17442242533e-11
R_2_110 n627 PAR_2_0_VDD075NNE 0.36016521471
R_3_110 PAR_3_1_VDD075NNE n628 2.32641290211
C_3_110 n628 PAR_2_0_VDD075NNE 8.11111324503e-11
L_4_110 PAR_3_1_VDD075NNE n629 1.91484113458e-09
R_4_110 n629 PAR_2_0_VDD075NNE 3.78760750172
R_5_110 PAR_3_1_VDD075NNE n630 10.1330413288
C_5_110 n630 PAR_2_0_VDD075NNE 1.27349563962e-10
L_6_110 PAR_3_1_VDD075NNE n631 3.36346291106e-07
R_6_110 n631 PAR_2_0_VDD075NNE 42.0534276916
G0_111 PAR_3_1_VDD075NNE PAR_3_0_VSS PAR_3_1_VDD075NNE PAR_3_0_VSS -2.2068282617
C0_111 PAR_3_1_VDD075NNE PAR_3_0_VSS 2.78863186149e-10
R_1_111 PAR_3_1_VDD075NNE n632 0.00494414994289
C_1_111 n632 PAR_3_0_VSS 3.37093745705e-09
R_2_111 PAR_3_1_VDD075NNE n633 0.0142406665179
C_2_111 n633 PAR_3_0_VSS 2.66180243198e-09
L_3_111 PAR_3_1_VDD075NNE n634 6.00466329581e-11
R_3_111 n634 PAR_3_0_VSS 0.453139020955
R_4_111 PAR_3_1_VDD075NNE n635 4.1962644843
C_4_111 n635 PAR_3_0_VSS 1.07143704233e-10
R_5_111 PAR_3_1_VDD075NNE n636 4.02819305843
C_5_111 n636 PAR_3_0_VSS 2.32676543771e-10
R_6_111 PAR_3_1_VDD075NNE n637 25.803504804
C_6_111 n637 PAR_3_0_VSS 3.85624470589e-10
R0_112 PAR_3_1_VDD075NNE PAR_3_0_VDD075NNE 0.00773794848576
C0_112 PAR_3_1_VDD075NNE PAR_3_0_VDD075NNE 2.66753018034e-10
L_1_112 PAR_3_1_VDD075NNE n638 3.70772703267e-13
R_1_112 n638 PAR_3_0_VDD075NNE 0.013748387564
L_2_112 PAR_3_1_VDD075NNE n639 4.1313728745e-12
R_2_112 n639 PAR_3_0_VDD075NNE 0.0788739226751
L_3_112 PAR_3_1_VDD075NNE n640 3.83886164674e-09
R_3_112 n640 PAR_3_0_VDD075NNE 14.9992466869
L_4_112 PAR_3_1_VDD075NNE n641 2.11022303227e-08
R_4_112 n641 PAR_3_0_VDD075NNE 31.3084839185
L_5_112 PAR_3_1_VDD075NNE n642 4.27301810144e-07
R_5_112 n642 PAR_3_0_VDD075NNE 204.391600882
L_6_112 PAR_3_1_VDD075NNE n643 0.00191092986457
R_6_112 n643 PAR_3_0_VDD075NNE 4725.51960665
G0_113 PAR_3_1_VDD075NNE PAR_0_1_VSS PAR_3_1_VDD075NNE PAR_0_1_VSS -2.32098636481
C0_113 PAR_3_1_VDD075NNE PAR_0_1_VSS 2.87849869804e-10
R_1_113 PAR_3_1_VDD075NNE n644 0.0503768457225
C_1_113 n644 PAR_0_1_VSS 3.08703375882e-10
L_2_113 PAR_3_1_VDD075NNE n645 7.21272023842e-11
R_2_113 n645 PAR_0_1_VSS 0.989133360886
L_3_113 PAR_3_1_VDD075NNE n646 2.26749571343e-10
R_3_113 n646 PAR_0_1_VSS 1.11896738407
L_4_113 PAR_3_1_VDD075NNE n647 1.43874675686e-09
R_4_113 n647 PAR_0_1_VSS 3.15939466345
L_5_113 PAR_3_1_VDD075NNE n648 1.30110520094e-08
R_5_113 n648 PAR_0_1_VSS 10.546359643
L_6_113 PAR_3_1_VDD075NNE n649 1.57708654524e-06
R_6_113 n649 PAR_0_1_VSS 200.663244148
G0_114 PAR_3_1_VDD075NNE PAR_0_1_VDD075NNE PAR_3_1_VDD075NNE PAR_0_1_VDD075NNE -8.70269052223
C0_114 PAR_3_1_VDD075NNE PAR_0_1_VDD075NNE 1.56164914724e-10
R_1_114 PAR_3_1_VDD075NNE n650 0.136940636879
C_1_114 n650 PAR_0_1_VDD075NNE 2.84894658713e-10
L_2_114 PAR_3_1_VDD075NNE n651 9.17038709411e-12
R_2_114 n651 PAR_0_1_VDD075NNE 0.130133370268
R_3_114 PAR_3_1_VDD075NNE n652 0.779576023789
C_3_114 n652 PAR_0_1_VDD075NNE 8.07484076063e-10
L_4_114 PAR_3_1_VDD075NNE n653 1.44216843594e-09
R_4_114 n653 PAR_0_1_VDD075NNE 0.981620538363
R_5_114 PAR_3_1_VDD075NNE n654 8.5100793002
C_5_114 n654 PAR_0_1_VDD075NNE 1.05879569863e-09
G0_115 PAR_3_1_VDD075NNE PAR_1_1_VSS PAR_3_1_VDD075NNE PAR_1_1_VSS -1.69537460268
C0_115 PAR_3_1_VDD075NNE PAR_1_1_VSS 2.89835307251e-10
R_1_115 PAR_3_1_VDD075NNE n655 0.0392808458546
C_1_115 n655 PAR_1_1_VSS 3.44580083659e-10
R_2_115 PAR_3_1_VDD075NNE n656 1.77134099541
C_2_115 n656 PAR_1_1_VSS 2.84572428832e-11
L_3_115 PAR_3_1_VDD075NNE n657 1.77575906857e-10
R_3_115 n657 PAR_1_1_VSS 0.961617931235
L_4_115 PAR_3_1_VDD075NNE n658 7.95557433368e-10
R_4_115 n658 PAR_1_1_VSS 1.96132036609
L_5_115 PAR_3_1_VDD075NNE n659 8.34880374201e-09
R_5_115 n659 PAR_1_1_VSS 7.2154424571
L_6_115 PAR_3_1_VDD075NNE n660 1.03544103179e-06
R_6_115 n660 PAR_1_1_VSS 142.68788917
G0_116 PAR_3_1_VDD075NNE PAR_1_1_VDD075NNE PAR_3_1_VDD075NNE PAR_1_1_VDD075NNE -8.59048777684
C0_116 PAR_3_1_VDD075NNE PAR_1_1_VDD075NNE 1.57821580377e-10
R_1_116 PAR_3_1_VDD075NNE n661 0.170385342611
C_1_116 n661 PAR_1_1_VDD075NNE 1.77366188832e-10
L_2_116 PAR_3_1_VDD075NNE n662 1.01864027252e-11
R_2_116 n662 PAR_1_1_VDD075NNE 0.147773140231
R_3_116 PAR_3_1_VDD075NNE n663 0.516543995757
C_3_116 n663 PAR_1_1_VDD075NNE 5.32786466934e-10
L_4_116 PAR_3_1_VDD075NNE n664 4.01735050506e-10
R_4_116 n664 PAR_1_1_VDD075NNE 0.59411759564
R_5_116 PAR_3_1_VDD075NNE n665 1.2730828745
C_5_116 n665 PAR_1_1_VDD075NNE 1.15393348716e-09
L_6_116 PAR_3_1_VDD075NNE n666 6.25189287195e-08
R_6_116 n666 PAR_1_1_VDD075NNE 7.16537906397
G0_117 PAR_3_1_VDD075NNE PAR_2_1_VSS PAR_3_1_VDD075NNE PAR_2_1_VSS -0.730187844224
C0_117 PAR_3_1_VDD075NNE PAR_2_1_VSS 2.36410632561e-10
R_1_117 PAR_3_1_VDD075NNE n667 0.0254416328402
C_1_117 n667 PAR_2_1_VSS 5.60950484631e-10
R_2_117 PAR_3_1_VDD075NNE n668 0.00962651471811
C_2_117 n668 PAR_2_1_VSS 3.85062727762e-09
R_3_117 PAR_3_1_VDD075NNE n669 2.18278026663
C_3_117 n669 PAR_2_1_VSS 6.25422756549e-11
L_4_117 PAR_3_1_VDD075NNE n670 6.941794282e-10
R_4_117 n670 PAR_2_1_VSS 1.74776430965
L_5_117 PAR_3_1_VDD075NNE n671 7.50904433017e-09
R_5_117 n671 PAR_2_1_VSS 6.64257494265
L_6_117 PAR_3_1_VDD075NNE n672 9.34265249724e-07
R_6_117 n672 PAR_2_1_VSS 133.613196264
R0_118 PAR_3_1_VDD075NNE PAR_2_1_VDD075NNE 0.00265920312619
C0_118 PAR_3_1_VDD075NNE PAR_2_1_VDD075NNE 1.55477058627e-10
L_1_118 PAR_3_1_VDD075NNE n673 2.98229106397e-13
R_1_118 n673 PAR_2_1_VDD075NNE 0.0137377665846
L_2_118 PAR_3_1_VDD075NNE n674 2.43816539475e-13
R_2_118 n674 PAR_2_1_VDD075NNE 0.00642451558774
L_3_118 PAR_3_1_VDD075NNE n675 1.03285088594e-10
R_3_118 n675 PAR_2_1_VDD075NNE 1.22255582694
L_4_118 PAR_3_1_VDD075NNE n676 1.82596572896e-08
R_4_118 n676 PAR_2_1_VDD075NNE 52.0960631203
L_5_118 PAR_3_1_VDD075NNE n677 1.23734296108e-07
R_5_118 n677 PAR_2_1_VDD075NNE 104.998212329
L_6_118 PAR_3_1_VDD075NNE n678 3.25394824791e-05
R_6_118 n678 PAR_2_1_VDD075NNE 2282.95056792
C0_119 PAR_3_1_VDD075NNE PAR_3_1_VSS 2.34959910533e-09
R_1_119 PAR_3_1_VDD075NNE n679 0.000328608821424
C_1_119 n679 PAR_3_1_VSS 5.6730924912e-08
R_2_119 PAR_3_1_VDD075NNE n680 0.000314125708188
C_2_119 n680 PAR_3_1_VSS 1.16417102973e-07
R_3_119 PAR_3_1_VDD075NNE n681 0.0863080106704
C_3_119 n681 PAR_3_1_VSS 1.35324400698e-09
R_4_119 PAR_3_1_VDD075NNE n682 0.665391716273
C_4_119 n682 PAR_3_1_VSS 5.81090385864e-10
R_5_119 PAR_3_1_VDD075NNE n683 26.9285319695
C_5_119 n683 PAR_3_1_VSS 4.37396596267e-10
G0_120 PAR_3_1_VDD075NNE PAR_0_0_VSS PAR_3_1_VDD075NNE PAR_0_0_VSS -0.988036366738
C0_120 PAR_3_1_VDD075NNE PAR_0_0_VSS 2.20900603745e-10
R_1_120 PAR_3_1_VDD075NNE n684 0.062838073768
C_1_120 n684 PAR_0_0_VSS 2.8209881287e-10
L_2_120 PAR_3_1_VDD075NNE n685 1.13423898683e-10
R_2_120 n685 PAR_0_0_VSS 1.05485546504
R_3_120 PAR_3_1_VDD075NNE n686 18.4601233761
C_3_120 n686 PAR_0_0_VSS 2.29808577505e-11
R_4_120 PAR_3_1_VDD075NNE n687 12.3068142802
C_4_120 n687 PAR_0_0_VSS 1.88068473246e-10
L_5_120 PAR_3_1_VDD075NNE n688 2.19935555509e-07
R_5_120 n688 PAR_0_0_VSS 24.9755268047
.ENDS

